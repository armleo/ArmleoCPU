
initial begin
	$dumpfile(`SIMRESULT);
	$dumpvars;
end
