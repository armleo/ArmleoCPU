////////////////////////////////////////////////////////////////////////////////
// 
// This file is part of ArmleoCPU.
// ArmleoCPU is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// ArmleoCPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with ArmleoCPU.  If not, see <https://www.gnu.org/licenses/>.
// 
// Copyright (C) 2016-2021, Arman Avetisyan, see COPYING file or LICENSE file
// SPDX-License-Identifier: GPL-3.0-or-later


// TODO: Add all undefs

`undef ACCESS_PACKED

`undef ARMLEOCPU_PAGE_METADATA_W
`undef ARMLEOCPU_PAGE_METADATA_VALID_BIT_NUM
`undef ARMLEOCPU_PAGE_METADATA_READ_BIT_NUM
`undef ARMLEOCPU_PAGE_METADATA_WRITE_BIT_NUM
`undef ARMLEOCPU_PAGE_METADATA_EXECUTE_BIT_NUM
`undef ARMLEOCPU_PAGE_METADATA_USER_BIT_NUM
`undef ARMLEOCPU_PAGE_METADATA_ACCESS_BIT_NUM
`undef ARMLEOCPU_PAGE_METADATA_DIRTY_BIT_NUM


`undef CACHE_RESPONSE_SUCCESS
`undef CACHE_RESPONSE_ACCESSFAULT
`undef CACHE_RESPONSE_PAGEFAULT
`undef CACHE_RESPONSE_MISSALIGNED
`undef CACHE_RESPONSE_UNKNOWNTYPE
`undef CACHE_RESPONSE_ATOMIC_FAIL


`undef AXI_BURST_INCR
`undef AXI_BURST_WRAP

`undef AXI_RESP_OKAY
`undef AXI_RESP_EXOKAY
`undef AXI_RESP_SLVERR
`undef AXI_RESP_DECERR

`undef CONNECT_AXI_BUS

`undef ARMLEOCPU_CSR_CMD_NONE
`undef ARMLEOCPU_CSR_CMD_READ
`undef ARMLEOCPU_CSR_CMD_WRITE
`undef ARMLEOCPU_CSR_CMD_READ_WRITE
`undef ARMLEOCPU_CSR_CMD_READ_SET
`undef ARMLEOCPU_CSR_CMD_READ_CLEAR
`undef ARMLEOCPU_CSR_CMD_MRET
`undef ARMLEOCPU_CSR_CMD_SRET
`undef ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN

`undef F2E_TYPE_WIDTH
`undef F2E_TYPE_INSTR
`undef F2E_TYPE_INTERRUPT_PENDING

`undef RD_ALU
`undef RD_CSR
`undef RD_DCACHE
`undef RD_LUI
`undef RD_AUIPC
`undef RD_PC_PLUS_4
`undef RD_MUL
`undef RD_MULH
`undef RD_DIV
`undef RD_REM
`undef RD_RS1
`undef RD_MINUS_ONE


`undef ARMLEOCPU_D2F_CMD_WIDTH
`undef ARMLEOCPU_D2F_CMD_FLUSH
`undef ARMLEOCPU_D2F_CMD_START_BRANCH
`undef ARMLEOCPU_D2F_CMD_NONE

`undef ARMLEOCPU_E2F_CMD_WIDTH
`undef ARMLEOCPU_E2F_CMD_FLUSH
`undef ARMLEOCPU_E2F_CMD_START_BRANCH
`undef ARMLEOCPU_E2F_CMD_NONE



`undef DEBUG_CMD_WIDTH
`undef DEBUG_CMD_NONE
`undef DEBUG_CMD_IFLUSH
`undef DEBUG_CMD_JUMP

`undef EXCEPTION_CODE_INTERRUPT
`undef INTERRUPT_CODE_SOFTWATE_INTERRUPT
`undef INTERRUPT_CODE_TIMER_INTERRUPT
`undef INTERRUPT_CODE_EXTERNAL_INTERRUPT

`undef EXCEPTION_CODE_SOFTWATE_INTERRUPT
`undef EXCEPTION_CODE_TIMER_INTERRUPT
`undef EXCEPTION_CODE_EXTERNAL_INTERRUPT

`undef EXCEPTION_CODE_INSTRUCTION_ADDRESS_MISSALIGNED
`undef EXCEPTION_CODE_INSTRUCTION_ACCESS_FAULT
`undef EXCEPTION_CODE_ILLEGAL_INSTRUCTION
`undef EXCEPTION_CODE_BREAKPOINT
`undef EXCEPTION_CODE_LOAD_ADDRESS_MISALIGNED
`undef EXCEPTION_CODE_LOAD_ACCESS_FAULT
`undef EXCEPTION_CODE_STORE_ADDRESS_MISALIGNED
`undef EXCEPTION_CODE_STORE_ACCESS_FAULT

`undef EXCEPTION_CODE_UCALL
`undef EXCEPTION_CODE_SCALL
`undef EXCEPTION_CODE_MCALL
`undef EXCEPTION_CODE_INSTRUCTION_PAGE_FAULT
`undef EXCEPTION_CODE_LOAD_PAGE_FAULT
`undef EXCEPTION_CODE_STORE_PAGE_FAULT


`undef INSTRUCTION_NOP


`undef OPCODE_LUI
`undef OPCODE_AUIPC
`undef OPCODE_JAL
`undef OPCODE_JALR
`undef OPCODE_BRANCH
`undef OPCODE_LOAD
`undef OPCODE_STORE
`undef OPCODE_OP_IMM
`undef OPCODE_OP
`undef OPCODE_FENCE
`undef OPCODE_SYSTEM

`undef ARMLEOCPU_PRIVILEGE_USER
`undef ARMLEOCPU_PRIVILEGE_USER_SV
`undef ARMLEOCPU_PRIVILEGE_SUPERVISOR
`undef ARMLEOCPU_PRIVILEGE_SUPERVISOR_SV
`undef ARMLEOCPU_PRIVILEGE_MACHINE


`undef TLB_CMD_NONE
`undef TLB_CMD_RESOLVE
`undef TLB_CMD_NEW_ENTRY
`undef TLB_CMD_INVALIDATE_ALL


`undef LOAD_BYTE
`undef LOAD_BYTE_UNSIGNED

`undef LOAD_HALF
`undef LOAD_HALF_UNSIGNED

`undef LOAD_WORD

`undef STORE_BYTE
`undef STORE_HALF
`undef STORE_WORD

`undef DEFINE_REG_REG_NXT
`undef DEFINE_CSR_REG
`undef DEFINE_CSR_OREG
`undef INIT_COMB_DEFAULT
`undef DEFINE_CSR_COMB_RO
`undef DEFINE_SCRATCH_CSR_REG_COMB
`undef DEFINE_ADDRESS_CSR_REG_COMB


`undef CHIP2CHIP_OPCODE_NONE
`undef CHIP2CHIP_OPCODE_READY
`undef CHIP2CHIP_OPCODE_WRITE

`default_nettype wire
