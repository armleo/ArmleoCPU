
// Here should be SDRAM Controller implementation
// But this implementation uses shared ADDR and DATA signals with multiple CS# signals
// This implementation is also compatible with io_share_unit