////////////////////////////////////////////////////////////////////////////////
// 
// This file is part of ArmleoCPU.
// ArmleoCPU is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// ArmleoCPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with ArmleoCPU.  If not, see <https://www.gnu.org/licenses/>.
// 
// Copyright (C) 2016-2021, Arman Avetisyan, see COPYING file or LICENSE file
// SPDX-License-Identifier: GPL-3.0-or-later
// 

/*
module armleocpu_decode (
// Fetch unit
    input      [31:0]       f2d_instr,
    input                   f2d_instr_valid,
    input      [31:0]       f2d_pc,
    input                   f2d_exc_start,
    input      [1:0]        f2d_exc_privilege,
    input      [31:0]       f2d_epc,
    input      [31:0]       f2d_cause,

    output reg              e2d_ready,
    output reg [`ARMLEOCPU_e2d_CMD_WIDTH-1:0]
                            e2d_cmd,
    output reg [31:0]       e2d_bubble_jump_target,
    output reg [31:0]       e2d_branchtarget,
);



endmodule*/
