`define ARMLEOCPU_E2F_CMD_WIDTH 2
`define ARMLEOCPU_E2F_CMD_BUBBLE_BRANCH (2'h3)
`define ARMLEOCPU_E2F_CMD_FLUSH (2'h2)
`define ARMLEOCPU_E2F_CMD_BRANCHTAKEN (2'h1)
`define ARMLEOCPU_E2F_CMD_IDLE (2'h0)