localparam EXCEPTION_CODE_INTERRUPT = 32'h8000_0000;
localparam EXCEPTION_CODE_SOFTWATE_INTERRUPT = 3 | EXCEPTION_CODE_INTERRUPT;
localparam EXCEPTION_CODE_TIMER_INTERRUPT = 7 | EXCEPTION_CODE_INTERRUPT;
localparam EXCEPTION_CODE_EXTERNAL_INTERRUPT = 11 | EXCEPTION_CODE_INTERRUPT;

localparam EXCEPTION_CODE_INSTRUCTION_ADDRESS_MISALIGNED = 0;
localparam EXCEPTION_CODE_INSTRUCTION_ACCESS_FAULT = 1;
localparam EXCEPTION_CODE_ILLEGAL_INSTRUCTION = 2;
localparam EXCEPTION_CODE_BREAKPOINT = 3;
localparam EXCEPTION_CODE_LOAD_ADDRESS_MISALIGNED = 4;
localparam EXCEPTION_CODE_LOAD_ACCESS_FAULT = 5;
localparam EXCEPTION_CODE_STORE_ADDRESS_MISALIGNED = 6;
localparam EXCEPTION_CODE_STORE_ACCESS_FAULT = 7;

// Calls from x privilege
localparam EXCEPTION_CODE_UCALL = 8;
localparam EXCEPTION_CODE_SCALL = 9;
localparam EXCEPTION_CODE_MCALL = 11;
localparam EXCEPTION_CODE_INSTRUCTION_PAGE_FAULT = 12;
localparam EXCEPTION_CODE_LOAD_PAGE_FAULT = 13;
localparam EXCEPTION_CODE_STORE_PAGE_FAULT = 15;
