////////////////////////////////////////////////////////////////////////////////
// 
// This file is part of ArmleoCPU.
// ArmleoCPU is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// ArmleoCPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with ArmleoCPU.  If not, see <https://www.gnu.org/licenses/>.
// 
// Copyright (C) 2016-2021, Arman Avetisyan, see COPYING file or LICENSE file
// SPDX-License-Identifier: GPL-3.0-or-later
// 
// Filename: armleocpu_csr.v
// Project:	ArmleoCPU
//
// Purpose:	CSR registers of ArmleoCPU,
//      also implements some interrupt related logic
//		
//
////////////////////////////////////////////////////////////////////////////////

`include "armleocpu_defines.vh"

`TIMESCALE_DEFINE

module armleocpu_csr(
    input clk,
    input rst_n,

    // Memory access level check registers
    // Used by multiple modules to calculate privilege level of current memory transaction
    output reg          csr_satp_mode,
    output reg [21:0]   csr_satp_ppn,

    output reg          csr_mstatus_mprv,
    output reg          csr_mstatus_mxr,
    output reg          csr_mstatus_sum,

    
    output reg [1:0]    csr_mstatus_mpp,
    output reg [1:0]    csr_mcurrent_privilege,

    // Trap registers
    // Used by execute to trap according instructions
    output reg          csr_mstatus_tsr,
    output reg          csr_mstatus_tw,
    output reg          csr_mstatus_tvm,

    // instret increment, generated by Execute unit
    input               instret_incr,


    // Interrupts logic, level sensitive
    input               irq_mtip_i, // Timer interrupt pending

    input               irq_meip_i,
    input               irq_seip_i,

    input               irq_mswi_i,
    input               irq_sswi_i,


    // Passed to fetch as "interrupt_pending" signal
    output reg          interrupt_pending_output,



    // Execute CSR commands and other related signals
    input      [3:0]    csr_cmd,

    output reg [31:0]   csr_next_pc,

    input      [11:0]   csr_address, // 12 bit address
    output reg          csr_invalid,
    // Shows that Invalid instruction should be generated

    output reg [31:0]   csr_to_rd, // Towards register
    input      [31:0]   csr_from_rs // From register
);



parameter MVENDORID = 32'h0A1AA1E0;
parameter MARCHID = 32'h1;
parameter MIMPID = 32'h1;
parameter MHARTID = 32'h0;



wire csr_write =    csr_cmd == `ARMLEOCPU_CSR_CMD_WRITE ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_WRITE ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_SET ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_CLEAR;

wire  csr_read =  csr_cmd == `ARMLEOCPU_CSR_CMD_READ ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_WRITE ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_SET ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_CLEAR;

`ifdef FORMAL_RULES
always @(posedge clk) begin
    assert(csr_read || csr_write || (csr_cmd == `ARMLEOCPU_CSR_CMD_NONE));
end
`endif

wire accesslevel_invalid = (csr_write || csr_read) && (csr_mcurrent_privilege < csr_address[9:8]);
wire write_invalid = (csr_write && (csr_address[11:10] == 2'b11));
reg csr_exists;

wire csr_invalid = accesslevel_invalid | write_invalid | csr_exists;

// holds read modify write operations first operand,
// because for mip, sip value used for RMW sequence is
// different from the value written to register

// See 3.1.9 Machine Interrupt Registers (mip and mie) in RISC-V Privileged spec

reg [31:0] rmw_before;
reg [31:0] rmw_after;


// TODO: Maybe make it REG instead of OREG because it's not connected to output
`DEFINE_CSR_OREG(32, csr_mtvec, 0)
`DEFINE_CSR_OREG(32, csr_stvec, 0)

`DEFINE_CSR_OREG(2, csr_mcurrent_privilege, 2'b11)
`DEFINE_CSR_OREG(1, csr_mstatus_tsr, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_tw, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_tvm, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_mxr, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_sum, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_mprv, 0)

`DEFINE_CSR_OREG(2, csr_mstatus_mpp, 0)
`DEFINE_CSR_REG(1, csr_mstatus_spp, 0)

`DEFINE_CSR_REG(1, csr_mstatus_mpie, 0)
`DEFINE_CSR_REG(1, csr_mstatus_spie, 0)

`DEFINE_CSR_REG(1, csr_mstatus_mie, 0)
`DEFINE_CSR_REG(1, csr_mstatus_sie, 0)

// MISA register logic below
`DEFINE_CSR_REG(1, csr_misa_atomic, 1)

`DEFINE_CSR_REG(32, csr_mscratch, 0)
`DEFINE_CSR_REG(32, csr_sscratch, 0)

`DEFINE_CSR_REG(32, csr_mepc, 0)
`DEFINE_CSR_REG(32, csr_sepc, 0)

`DEFINE_CSR_REG(32, csr_mcause, 0)
`DEFINE_CSR_REG(32, csr_scause, 0)

`DEFINE_CSR_REG(32, csr_mtval, 0)
`DEFINE_CSR_REG(32, csr_stval, 0)

`DEFINE_CSR_REG(32, csr_cycle, 0)
`DEFINE_CSR_REG(32, csr_cycleh, 0)

`DEFINE_CSR_REG(32, csr_instret, 0)
`DEFINE_CSR_REG(32, csr_instreth, 0)

`DEFINE_CSR_OREG(22, csr_satp_ppn, 0)
`DEFINE_CSR_OREG(1, csr_satp_mode, 0)

`DEFINE_CSR_OREG(16, csr_medeleg, 0)
`DEFINE_CSR_OREG(12, csr_mideleg, 0)

wire csr_mideleg_external_interrupt = csr_mideleg[9];
wire csr_mideleg_timer_interrupt = csr_mideleg[5];
wire csr_mideleg_software_interrupt = csr_mideleg[1];

`DEFINE_CSR_REG(1, csr_mie_meie, 0)
// 11th bit, active and read/writeable when no mideleg
`DEFINE_CSR_REG(1, csr_mie_seie, 0)
// 9th bit, active and read/writeable when mideleg

`DEFINE_CSR_REG(1, csr_mie_mtie, 0)
// 7th bit, active and read/writeable when no mideleg
`DEFINE_CSR_REG(1, csr_mie_stie, 0)
// 5th bit, active and read/writeable when mideleg

`DEFINE_CSR_REG(1, csr_mie_msie, 0)
// 3th bit, active and read/writeable when no mideleg

`DEFINE_CSR_REG(1, csr_mie_ssie, 0)
// 1th bit, active and read/writeable when mideleg

`DEFINE_CSR_REG(1, csr_mip_seip, 0)
// 9th bit, read/write if mideleg, else zero
// when read seip is logical or of this bit and external signal
// when rmw then seip is this bit

`DEFINE_CSR_REG(1, csr_mip_stip, 0)
// 5th bit, read/write if mideleg, else zero
`DEFINE_CSR_REG(1, csr_mip_ssip, 0)
// 1th bit, read/write if mideleg, else zero


wire [31:0] csr_misa = {
    2'b01, // MXLEN = 32, only valid value
    4'b0000, // Reserved
    1'b0, // Z
    1'b0, // Y
    1'b0, // X
    1'b0, // W
    1'b0, // V
    1'b1, // U - User mode, present
    1'b0, // T
    1'b1, // S - Supervisor mode, present
    1'b0, // R
    1'b0, // Q
    1'b0, // P
    1'b0, // O
    1'b0, // N
    1'b1, // M - Multiply/Divide, Present
    1'b0, // L
    1'b0, // K
    1'b0, // J
    1'b1, // I - RV32I
    1'b0, // H
    1'b0, // G
    1'b0, // F
    1'b0, // E
    1'b0, // D
    1'b0, // C
    1'b0, // B
    csr_misa_atomic  // A
};


// This signal is calculated SIE
// It is calculated because this signal is low
// To block supervisor level interrupts in machine mode
reg supervisor_user_calculated_sie;


always @* begin
    rmw_after = csr_from_rs;
    if(csr_cmd == `ARMLEOCPU_CSR_CMD_READ_WRITE || csr_cmd == `ARMLEOCPU_CSR_CMD_WRITE)
        rmw_after = csr_from_rs;
    else if(csr_cmd == `ARMLEOCPU_CSR_CMD_READ_SET)
        rmw_after = rmw_before | csr_from_rs;
    else if(csr_cmd == `ARMLEOCPU_CSR_CMD_READ_CLEAR)
        rmw_after = rmw_before & ~csr_from_rs;
    // We don't care about this signal in read only operations
    // Because no write is done for this operations
end


// TODO: output next_pc


always @* begin

    csr_exists = 0;
    csr_to_rd = 0;

    // TODO: Add all default values for macros above
    

    {csr_instreth_nxt, csr_instret_nxt} = {csr_instreth, csr_instret} + instret_incr;
    {csr_cycleh_nxt, csr_cycle_nxt} = {csr_cycleh, csr_cycle} + 1;
end

endmodule

`include "armleocpu_undef.vh"
