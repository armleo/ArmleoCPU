////////////////////////////////////////////////////////////////////////////////
// 
// This file is part of ArmleoCPU.
// ArmleoCPU is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// ArmleoCPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with ArmleoCPU.  If not, see <https://www.gnu.org/licenses/>.
// 
// Copyright (C) 2016-2021, Arman Avetisyan, see COPYING file or LICENSE file
// SPDX-License-Identifier: GPL-3.0-or-later
// 
// Note: ADDR_WIDTH is fixed to 32 bits.
//      All unused bits can be assigned to zero
//      
// Implementation details:
//      AXI bus is registered (bus_upstream_axi_* <-> upstream_axi_*)
//      An clock is generated on the output.
//      clk signal of this module is divided by two and connected to
//      clk_enable signal. This signal is used by logic below to control
//      IO signals.
//      As clk can be running at higher or same frequency than
//      data clock is used by device.
//      Output clock is generated by
//      
//      
//      When bus changes direction io_oe is asserted/deasserted,
//      then both sides wait single cycle.
//      And then starting to accept the data.
//      It is possible for bus to be in Hi-Z state,
//      but both OE's assertion is impossible.
//      
//      For each AXI write request we write all write data and aw* data
//      into temporary storage. Then owned_by_bus is reset.
//      Same is done for AXI read requests, except no write data is set
//      
//      Why store AXI request in buffer anyway?
//      AXI Does not guarantee that Write data will be provided every cycle
//      This makes possible the scenario when write data valid is
//      deasserted, causing no data to be available.
//      So instead of making it a requirement we just buffer it.
//      
//      
//      If any buffer has owned_by_bus reset then following logic is executed
//      1. CSN is asserted (CSN=0 is because its inverted) by host.
//      2. Bus logic starts transmission of packet. (up to 8 + 16*32 cycles)
//      3. Bus logic de-asserts OE for two cycles. Device asserts OE
//      4. Host waits for response packet start
//          Note:(While bus is idle all bits are low)
//      5. Device sends response when ready
//      6. Device drives Hi-Z on the bus
//      7. Host waits two cycles and asserts bus with all-zero,
//          CSN is asserted high.
//      
//      Multiple types of packets are possible
//      WRITE/READ/SYNC
//      Sync is used by host to poll IRQ bit
//      Write is write request
//      Read is read request
//      Each packet structure is provided in code below
//      
////////////////////////////////////////////////////////////////////////////////

`include "armleocpu_defines.vh"

`TIMESCALE_DEFINE

module armleocpu_chip2chip_host(
    clk, rst_n,

    bus_upstream_axi_awvalid, bus_upstream_axi_awready, bus_upstream_axi_awaddr, bus_upstream_axi_awlen, bus_upstream_axi_awburst, bus_upstream_axi_awsize,
    bus_upstream_axi_wvalid, bus_upstream_axi_wready, bus_upstream_axi_wdata, bus_upstream_axi_wstrb, bus_upstream_axi_wlast,
    bus_upstream_axi_bvalid, bus_upstream_axi_bready, bus_upstream_axi_bresp,

    bus_upstream_axi_arvalid, bus_upstream_axi_arready, bus_upstream_axi_araddr, bus_upstream_axi_arlen, bus_upstream_axi_arsize, bus_upstream_axi_arburst,
    bus_upstream_axi_rvalid, bus_upstream_axi_rready, bus_upstream_axi_rresp, bus_upstream_axi_rlast, bus_upstream_axi_rdata,

    bus_upstream_irq,

    // TODO: Add signals
);

parameter ID_WIDTH = 4;
localparam ADDR_WIDTH = 32;
localparam DATA_WIDTH = 32;
localparam DATA_STROBES = DATA_WIDTH/8;

input                   clk;
input                   rst_n;

output reg                      bus_upstream_irq;

input wire                      bus_upstream_axi_awvalid;
output wire                     bus_upstream_axi_awready;
input wire  [ADDR_WIDTH-1:0]    bus_upstream_axi_awaddr;
input wire  [7:0]               bus_upstream_axi_awlen;
input wire  [SIZE_WIDTH-1:0]    bus_upstream_axi_awsize;
input wire  [1:0]               bus_upstream_axi_awburst;
input wire                      bus_upstream_axi_awlock;
input wire  [ID_WIDTH-1:0]      bus_upstream_axi_awid;
input wire  [2:0]               bus_upstream_axi_awprot;

// AXI W Bus
input wire                      bus_upstream_axi_wvalid;
output wire                     bus_upstream_axi_wready;
input wire  [DATA_WIDTH-1:0]    bus_upstream_axi_wdata;
input wire  [DATA_STROBES-1:0]  bus_upstream_axi_wstrb;
input wire                      bus_upstream_axi_wlast;

// AXI B Bus
output wire                     bus_upstream_axi_bvalid;
input wire                      bus_upstream_axi_bready;
output wire [1:0]               bus_upstream_axi_bresp;
output wire [ID_WIDTH-1:0]      bus_upstream_axi_bid;

input wire                      bus_upstream_axi_arvalid;
output wire                     bus_upstream_axi_arready;
input wire  [ADDR_WIDTH-1:0]    bus_upstream_axi_araddr;
input wire  [7:0]               bus_upstream_axi_arlen;
input wire  [SIZE_WIDTH-1:0]    bus_upstream_axi_arsize;
input wire  [1:0]               bus_upstream_axi_arburst;
input wire  [ID_WIDTH-1:0]      bus_upstream_axi_arid;
input wire                      bus_upstream_axi_arlock;
input wire  [2:0]               bus_upstream_axi_arprot;

output wire                     bus_upstream_axi_rvalid;
input  wire                     bus_upstream_axi_rready;
output wire [1:0]               bus_upstream_axi_rresp;
output wire                     bus_upstream_axi_rlast;
output wire [DATA_WIDTH-1:0]    bus_upstream_axi_rdata;
output wire [ID_WIDTH-1:0]      bus_upstream_axi_rid;

// TODO: Add ctrl AXI4 bus.
// This ctrl bus is used to control frequency.

output reg  [0:0]               io_csn;
input wire  [7:0]               io_datain;
output reg  [7:0]               io_dataout;
output reg                      io_oe;
output reg                      io_clk_out;



armleocpu_axi_register_slice #(
    .ADDR_WIDTH(ADDR_WIDTH), // Fixed
    .ID_WIDTH(ID_WIDTH), // Configurable
    .DATA_WIDTH(DATA_WIDTH) // Fixed
) slice(
    .clk                (clk),
    .rst_n              (rst_n),

    `CONNECT_AXI_BUS(upstream_axi_, bus_upstream_axi_)
    .upstream_axi_arlock           (io_upstream_arlock),
    .upstream_axi_awlock           (io_upstream_awlock),

    `CONNECT_AXI_BUS(downstream_axi_, upstream_axi_), 
    .downstream_axi_arlock         (upstream_axi_arlock),
    .downstream_axi_awlock         (upstream_axi_awlock),
);



reg [4:0] address;

armleocpu_mem_1rw #(
    .ELEMENTS_W(5), // at least (8 + 16) x 32 -> rounded up 32 x 32
    .WIDTH(DATA_WIDTH),
) buffer0 (
    .clk        (clk),

    .address    (address),

    .read       (read),
    .readdata   (readdata),

    .write      (write),
    .writedata  (writedata)
);



always @* begin

    state_nxt = state;
    address = 0;
    write = 0;
    read = 0;
    writedata = 0;

    upstream_axi_awready = 0;
    upstream_axi_wready = 0;
    upstream_axi_bvalid = 0;
    upstream_axi_arready = 0;
    upstream_axi_rvalid = 0;

    currently_writing_nxt = currently_writing;

    case(state)
        STATE_IDLE: begin
            address = 0;
            if(upstream_axi_awvalid) begin
                writedata = {, OPCODE_WRITE};
                write = 1;
                currently_writing_nxt = 1;
                `ifdef DEBUG_CHIP2CHIP
                assume(upstream_axi_awlen < 16); // Make sure no bigger than 64 bytes per burst
                `endif
            end else if(upstream_axi_arvalid) begin
                writedata = OPCODE_READ;
                write = 1;
                currently_writing_nxt = 0;
                `ifdef DEBUG_CHIP2CHIP
                assume(upstream_axi_arlen < 16); // Make sure no bigger than 64 bytes per burst
                `endif
            end
        end
        
        STATE_WRITE0: begin
            write = 1;
            address = 1;
            if(currently_writing) begin // AW
                writedata = {
                    upstream_axi_awaddr, // 32 bits
                };
            end else begin // AR
                writedata = {
                    upstream_axi_araddr
                };
            end

            state_nxt = STATE_WRITE1;
        end
        STATE_WRITE1: begin
            write = 1;
            
            address = 2;
            if(currently_writing) begin
                writedata = {
                    upstream_axi_awid,   // ID_WIDTH
                    upstream_axi_awlen,  // 8
                    upstream_axi_awsize, // 3
                    upstream_axi_awburst,// 2
                    upstream_axi_awlock, // 1
                    upstream_axi_awprot  // 3
                };
            end else begin
                writedata = {
                    upstream_axi_awid,   // ID_WIDTH
                    upstream_axi_awlen,  // 8
                    upstream_axi_awsize, // 3
                    upstream_axi_awburst,// 2
                    upstream_axi_awlock, // 1
                    upstream_axi_awprot  // 3
                };
            end


            state_nxt = STATE_WRITE_DATA;

            len_nxt = len;
        end
        STATE_WRITE_DATA: begin
            
            if()
            counter_nxt = 2 + len;
            state_nxt = STATE_TX;
            initial_cycle_nxt = 1;
        end
        STATE_TX: begin
            io_csn = 0;
            
            read = 1;
            initial_cycle_nxt = 0;
            if(initial_cycle) begin
                
            end else if(counter != 0) begin

            else begin

            end
            
            state_nxt = STATE_RX;
        end
        STATE_RX: begin

            state_nxt = STATE_IDLE;
        end
    endcase
end




endmodule


`include "armleocpu_undef.vh"
