parameter RESET_VECTOR = 32'h0000_0000;