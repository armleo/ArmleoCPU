`define CACHE_RESPONSE_IDLE 4'd0
`define CACHE_RESPONSE_WAIT 4'd1
`define CACHE_RESPONSE_DONE 4'd2
`define CACHE_RESPONSE_ACCESSFAULT 4'd3
`define CACHE_RESPONSE_PAGEFAULT 4'd4
`define CACHE_RESPONSE_MISSALIGNED 4'd5
`define CACHE_RESPONSE_UNKNOWNTYPE 4'd6

`define CACHE_CMD_NONE 4'd0
`define CACHE_CMD_EXECUTE 4'd1
`define CACHE_CMD_LOAD 4'd2
`define CACHE_CMD_STORE 4'd3
`define CACHE_CMD_FLUSH_ALL 4'd4


