`define ARMLEOBUS_CMD_NONE 3'd0
`define ARMLEOBUS_CMD_READ 3'd1
`define ARMLEOBUS_CMD_WRITE 3'd2

`define CACHE_CMD_NONE 3'd0
`define CACHE_CMD_EXECUTE 3'd1
`define CACHE_CMD_LOAD 3'd2
`define CACHE_CMD_STORE 3'd3
