////////////////////////////////////////////////////////////////////////////////
// 
// This file is part of ArmleoCPU.
// ArmleoCPU is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
// 
// ArmleoCPU is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with ArmleoCPU.  If not, see <https://www.gnu.org/licenses/>.
// 
// Copyright (C) 2016-2021, Arman Avetisyan, see COPYING file or LICENSE file
// SPDX-License-Identifier: GPL-3.0-or-later
// 
// Filename: armleocpu_csr.v
// Project:	ArmleoCPU
//
// Purpose:	CSR registers of ArmleoCPU,
//      also implements some interrupt related logic
//		
//
////////////////////////////////////////////////////////////////////////////////

`include "armleocpu_defines.vh"

`TIMESCALE_DEFINE

module armleocpu_csr(
    input wire clk,
    input wire rst_n,

    // Memory access level check registers
    // Used by multiple modules to calculate privilege level of current memory transaction
    output reg          csr_satp_mode,
    output reg [21:0]   csr_satp_ppn,

    output reg          csr_mstatus_mprv,
    output reg          csr_mstatus_mxr,
    output reg          csr_mstatus_sum,

    
    output reg [1:0]    csr_mstatus_mpp,
    output reg [1:0]    csr_mcurrent_privilege,

    // Trap registers
    // Used by execute to trap according instructions
    output reg          csr_mstatus_tsr,
    output reg          csr_mstatus_tw,
    output reg          csr_mstatus_tvm,

    // instret increment, generated by Execute unit
    // Assumed sync to clk
    input wire          instret_incr,


    // Interrupts logic, level sensitive
    input wire          irq_mtip_i, // Timer interrupt pending
    input wire          irq_stip_i, // Might as well keep it, because logic is implemented anyway
    // If stip is not implemented, just tie it to zero

    input wire          irq_meip_i, // External interrupt pending
    input wire          irq_seip_i,

    input wire          irq_msip_i, // Software interrupt pending
    input wire          irq_ssip_i,


    // Passed to fetch as "interrupt_pending" signal
    // Fetch when starts new fetch and detects this signal asserted
    // then no fetch is issued and "interrupt pending" f2d packet is
    // passed to decode stage.
    // Decode stage then passes it to Execute stage
    // Then execute stage issues csr_cmd INTERRUPT_BEGIN
    output reg          interrupt_pending_output,




    // Note: outputs are changed only after cycle that csr_cmd retires
    //      This means that before jumping to csr_next_pc has
    //      to wait for CSR_CMD to retire.
    //      
    //      Also worth mentioning that execute module should not rely
    //      on any of CSR outputs until first instruction from csr_next_pc.
    //
    //      Implementations must ensure that once CSR_CMD is retired
    //      None of CSR outputs influence the execute unit's outcome
    //      
    //      Example: SRET is executed. CSR_CMD is signaled and csr_next_pc is registered
    //      Problem arises in case that for example execute relies on csr_mcurrent_privilege
    //      As on second cycle this is now set to value of PP causing pagefault
    //      Which is an issue. Instead Execute implementation should raise a flag
    //      When this flag is raised then execute just does e2d command
    //      Ignoring all CSR outputs

    // Execute CSR commands and other related signals
    input wire [3:0]    csr_cmd,

    
    // Used to signal execute where to continue execution from
    output reg [31:0]   csr_next_pc,
    input wire [31:0]   csr_exc_epc,
    input wire [31:0]   csr_exc_cause,

    input wire [11:0]   csr_address, // 12 bit address
    output wire         csr_cmd_error,
    // Shows that Invalid instruction should be generated

    output reg [31:0]   csr_to_rd, // Towards register
    input wire [31:0]   csr_from_rs // From register
);



parameter [31:0] MVENDORID = 32'h0A1AA1E0;
parameter [31:0] MARCHID = 32'h1;
parameter [31:0] MIMPID = 32'h1;
parameter [31:0] MHARTID = 32'h0;
parameter [31:0] MCONFIGPTR = 32'h100;


wire csr_write =    csr_cmd == `ARMLEOCPU_CSR_CMD_WRITE ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_WRITE ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_SET ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_CLEAR;

wire  csr_read =  csr_cmd == `ARMLEOCPU_CSR_CMD_READ ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_WRITE ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_SET ||
                    csr_cmd == `ARMLEOCPU_CSR_CMD_READ_CLEAR;

`ifdef FORMAL_RULES
always @(posedge clk) begin
    assert(
        csr_read || csr_write
        || (csr_cmd == `ARMLEOCPU_CSR_CMD_NONE)
        || (csr_cmd == `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN)
        || (csr_cmd == `ARMLEOCPU_CSR_CMD_MRET)
        || (csr_cmd == `ARMLEOCPU_CSR_CMD_SRET)
    );
end
`endif

wire accesslevel_invalid = (csr_write || csr_read) && (csr_mcurrent_privilege < csr_address[9:8]);
wire write_invalid = (csr_write && (csr_address[11:10] == 2'b11));
reg csr_exists;


wire csr_invalid = (csr_read || csr_write) && (accesslevel_invalid | write_invalid | !csr_exists);

reg csr_cmd_exc_int_error;

assign csr_cmd_error = csr_invalid | csr_cmd_exc_int_error;




// holds read modify write operations first operand,
// because for mip, sip value used for RMW sequence is
// different from the value written to register

// See 3.1.9 Machine Interrupt Registers (mip and mie) in RISC-V Privileged spec

// verilator coverage_off
reg [31:0] rmw_before;
reg [31:0] rmw_after;


`DEFINE_CSR_REG(32, csr_mtvec, 0)
`DEFINE_CSR_REG(32, csr_stvec, 0)

`DEFINE_CSR_OREG(2, csr_mcurrent_privilege, 2'b11)
`DEFINE_CSR_OREG(1, csr_mstatus_tsr, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_tw, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_tvm, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_mxr, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_sum, 0)
`DEFINE_CSR_OREG(1, csr_mstatus_mprv, 0)

`DEFINE_CSR_OREG(2, csr_mstatus_mpp, 0)
`DEFINE_CSR_REG(1, csr_mstatus_spp, 0)

`DEFINE_CSR_REG(1, csr_mstatus_mpie, 0)
`DEFINE_CSR_REG(1, csr_mstatus_spie, 0)

`DEFINE_CSR_REG(1, csr_mstatus_mie, 0)
`DEFINE_CSR_REG(1, csr_mstatus_sie, 0)

`DEFINE_CSR_REG(32, csr_mscratch, 0)
`DEFINE_CSR_REG(32, csr_sscratch, 0)

`DEFINE_CSR_REG(32, csr_mepc, 0)
`DEFINE_CSR_REG(32, csr_sepc, 0)

`DEFINE_CSR_REG(32, csr_mcause, 0)
`DEFINE_CSR_REG(32, csr_scause, 0)

// MTVAL is allowed to be hardwired to zero, if never written
// STVAL CANT BE hardwired to zero
`DEFINE_CSR_REG(32, csr_stval, 0)

`DEFINE_CSR_REG(32, csr_cycle, 0)
`DEFINE_CSR_REG(32, csr_cycleh, 0)

`DEFINE_CSR_REG(32, csr_instret, 0)
`DEFINE_CSR_REG(32, csr_instreth, 0)

`DEFINE_CSR_OREG(22, csr_satp_ppn, 0)
`DEFINE_CSR_OREG(1, csr_satp_mode, 0)


`DEFINE_CSR_REG(1, csr_mie_meie, 0)
// 11th bit, active and read/writeable when no mideleg
`DEFINE_CSR_REG(1, csr_mie_seie, 0)
// 9th bit, active and read/writeable when mideleg

`DEFINE_CSR_REG(1, csr_mie_mtie, 0)
// 7th bit, active and read/writeable when no mideleg
`DEFINE_CSR_REG(1, csr_mie_stie, 0)
// 5th bit, active and read/writeable when mideleg

`DEFINE_CSR_REG(1, csr_mie_msie, 0)
// 3th bit, active and read/writeable when no mideleg

`DEFINE_CSR_REG(1, csr_mie_ssie, 0)
// 1th bit, active and read/writeable when mideleg



`DEFINE_CSR_REG(1, csr_mip_seip, 0)
// 9th bit, read/write if mideleg, else zero
// when read seip is logical or of this bit and external signal
// when rmw then seip is this bit
// csr_mip_meip does not exist because is read only


`DEFINE_CSR_REG(1, csr_mip_stip, 0)
// 5th bit, read/write if mideleg, else zero
`DEFINE_CSR_REG(1, csr_mip_ssip, 0)
// 1th bit, read/write if mideleg, else zero

wire [31:0] csr_misa = {
    2'b01, // MXLEN = 32, only valid value
    4'b0000, // Reserved
    1'b0, // Z
    1'b0, // Y
    1'b0, // X
    1'b0, // W
    1'b0, // V
    1'b1, // U - User mode, present
    1'b0, // T
    1'b1, // S - Supervisor mode, present
    1'b0, // R
    1'b0, // Q
    1'b0, // P
    1'b0, // O
    1'b0, // N
    1'b1, // M - Multiply/Divide, Present
    1'b0, // L
    1'b0, // K
    1'b0, // J
    1'b1, // I - RV32I
    1'b0, // H
    1'b0, // G
    1'b0, // F
    1'b0, // E
    1'b0, // D
    1'b0, // C
    1'b0, // B
    1'b1  // A
};
// verilator coverage_on

// This signal is calculated SIE
// It is calculated because this signal is low
// To block supervisor level interrupts in machine mode
reg supervisor_user_calculated_sie;
reg machine_calculated_mie;

reg irq_calculated_meie;
reg irq_calculated_mtie;
reg irq_calculated_msie;

reg irq_calculated_seie;
reg irq_calculated_stie;
reg irq_calculated_ssie;

// pending
reg irq_calculated_meip;
reg irq_calculated_mtip;
reg irq_calculated_msip;

reg irq_calculated_seip;
reg irq_calculated_stip;
reg irq_calculated_ssip;

// verilator coverage_off
always @* begin
    rmw_after = csr_from_rs;
    // verilator coverage_on
    if(csr_cmd == `ARMLEOCPU_CSR_CMD_READ_WRITE || csr_cmd == `ARMLEOCPU_CSR_CMD_WRITE)
        rmw_after = csr_from_rs;
    else if(csr_cmd == `ARMLEOCPU_CSR_CMD_READ_SET)
        rmw_after = rmw_before | csr_from_rs;
    else if(csr_cmd == `ARMLEOCPU_CSR_CMD_READ_CLEAR)
        rmw_after = rmw_before & ~csr_from_rs;
    // We don't care about this signal in read only operations
    // Because no write is done for this operations
end

wire csr_mcurrent_privilege_machine = csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_MACHINE;
wire csr_mcurrent_privilege_supervisor = csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_SUPERVISOR;
wire csr_mcurrent_privilege_machine_supervisor = csr_mcurrent_privilege_machine | csr_mcurrent_privilege_supervisor;

// verilator coverage_off
always @* begin

    csr_exists = 0;
    csr_to_rd = 0;

    rmw_before = 0;
    csr_next_pc = csr_mtvec;

    // Note: csr_invalid is only check for privilege
    // and write allowing

    // Only signal assigned to error return is
    // csr_exists, which is set when we are not able to find
    // csr for that specific address
    
    `INIT_COMB_DEFAULT(csr_mtvec)
    `INIT_COMB_DEFAULT(csr_stvec)
    `INIT_COMB_DEFAULT(csr_mcurrent_privilege)

    // Note: sstatus is limited representation of mstatus
    // so no separate set of registers are required
    // to implement them
    
    `INIT_COMB_DEFAULT(csr_mstatus_tsr)
    `INIT_COMB_DEFAULT(csr_mstatus_tw)
    `INIT_COMB_DEFAULT(csr_mstatus_tvm)
    `INIT_COMB_DEFAULT(csr_mstatus_mxr)
    `INIT_COMB_DEFAULT(csr_mstatus_sum)
    `INIT_COMB_DEFAULT(csr_mstatus_mprv)
    `INIT_COMB_DEFAULT(csr_mstatus_mpp)
    `INIT_COMB_DEFAULT(csr_mstatus_spp)
    `INIT_COMB_DEFAULT(csr_mstatus_mpie)
    `INIT_COMB_DEFAULT(csr_mstatus_spie)
    `INIT_COMB_DEFAULT(csr_mstatus_mie)
    `INIT_COMB_DEFAULT(csr_mstatus_sie)

    `INIT_COMB_DEFAULT(csr_mscratch)
    `INIT_COMB_DEFAULT(csr_sscratch)
    `INIT_COMB_DEFAULT(csr_mepc)
    `INIT_COMB_DEFAULT(csr_sepc)
    `INIT_COMB_DEFAULT(csr_mcause)
    `INIT_COMB_DEFAULT(csr_scause)
    `INIT_COMB_DEFAULT(csr_stval)

    // cycle and instret skipped, assigned in logic below

    `INIT_COMB_DEFAULT(csr_satp_ppn)
    `INIT_COMB_DEFAULT(csr_satp_mode)

    `INIT_COMB_DEFAULT(csr_mie_meie)
    `INIT_COMB_DEFAULT(csr_mie_seie)

    `INIT_COMB_DEFAULT(csr_mie_mtie)
    `INIT_COMB_DEFAULT(csr_mie_stie)

    `INIT_COMB_DEFAULT(csr_mie_msie)
    `INIT_COMB_DEFAULT(csr_mie_ssie)

    // csr_mip_meip does not exist because is read only
    `INIT_COMB_DEFAULT(csr_mip_seip)

    `INIT_COMB_DEFAULT(csr_mip_stip)
    `INIT_COMB_DEFAULT(csr_mip_ssip)

    // TODO: Add all default values for macros above
    
    // Interrupt handling related signals
    
    

    // verilator lint_off WIDTH
    {csr_instreth_nxt, csr_instret_nxt} = {csr_instreth, csr_instret} + instret_incr;
    // verilator lint_on WIDTH
    {csr_cycleh_nxt, csr_cycle_nxt} = {csr_cycleh, csr_cycle} + 1;
    
    

    // Interrupt enabled/disabled section
    // Logic below is as following:
    // Calculated M*IE signals are as follows
    //  if machine mode then use MIE and M*IE
    //  if supervisor/user mode then ignore MIE and use M*IE only
    // Calculated S*IE signals are as follows
    //  if supervisor mode then use S*IE and SIE
    //  if user mode then only use S*IE
    //  if machine just disable

    machine_calculated_mie =
        (
            (csr_mcurrent_privilege_machine)
            & csr_mstatus_mie
        ) | (!csr_mcurrent_privilege_machine);

    irq_calculated_meie = machine_calculated_mie & csr_mie_meie;
    irq_calculated_mtie = machine_calculated_mie & csr_mie_mtie;
    irq_calculated_msie = machine_calculated_mie & csr_mie_msie;


    supervisor_user_calculated_sie =
        (
            (csr_mcurrent_privilege_supervisor)
            & csr_mstatus_sie
        ) | (csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_USER);

    irq_calculated_seie = supervisor_user_calculated_sie & csr_mie_seie;
    irq_calculated_stie = supervisor_user_calculated_sie & csr_mie_stie;
    irq_calculated_ssie = supervisor_user_calculated_sie & csr_mie_ssie;

    
    irq_calculated_meip = irq_meip_i;
    irq_calculated_mtip = irq_mtip_i;
    irq_calculated_msip = irq_msip_i;

    irq_calculated_seip = irq_seip_i | csr_mip_seip;
    irq_calculated_stip = irq_stip_i | csr_mip_stip;
    irq_calculated_ssip = irq_ssip_i | csr_mip_ssip;

    interrupt_pending_output = 
        (irq_calculated_meip & irq_calculated_meie) |
        (irq_calculated_mtip & irq_calculated_mtie) |
        (irq_calculated_msip & irq_calculated_msie) |
        (irq_calculated_seip & irq_calculated_seie) |
        (irq_calculated_stip & irq_calculated_stie) |
        (irq_calculated_ssip & irq_calculated_ssie);


    csr_cmd_exc_int_error = 1;

    // verilator coverage_on

    if(csr_cmd == `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN) begin
        // Note: Order matters, checkout the interrupt priority in RISC-V Privileged Manual
        if(irq_calculated_meip & irq_calculated_meie) begin // MEI
            csr_mcause_nxt = `EXCEPTION_CODE_MACHINE_EXTERNAL_INTERRUPT; // Calculated by the CSR
            csr_cmd_exc_int_error = 0;
        end else if(irq_calculated_msip & irq_calculated_msie) begin // MSI
            csr_mcause_nxt = `EXCEPTION_CODE_MACHINE_SOFTWATE_INTERRUPT; // Calculated by the CSR
            csr_cmd_exc_int_error = 0;
        end else if(irq_calculated_mtip & irq_calculated_mtie) begin // MTI
            csr_mcause_nxt = `EXCEPTION_CODE_MACHINE_TIMER_INTERRUPT; // Calculated by the CSR
            csr_cmd_exc_int_error = 0;
        end else if(irq_calculated_seip & irq_calculated_seie) begin // SEI
            csr_mcause_nxt = `EXCEPTION_CODE_SUPERVISOR_EXTERNAL_INTERRUPT; // Calculated by the CSR
            csr_cmd_exc_int_error = 0;
        end else if(irq_calculated_ssip & irq_calculated_ssie) begin // SSI
            csr_mcause_nxt = `EXCEPTION_CODE_SUPERVISOR_SOFTWATE_INTERRUPT; // Calculated by the CSR
            csr_cmd_exc_int_error = 0;
        end else if(irq_calculated_stip & irq_calculated_stie) begin // STI
            csr_mcause_nxt = `EXCEPTION_CODE_SUPERVISOR_TIMER_INTERRUPT; // Calculated by the CSR
            csr_cmd_exc_int_error = 0;
        end else begin
            csr_cmd_exc_int_error = 1;
        end

        if(!csr_cmd_exc_int_error) begin
            csr_mstatus_mpie_nxt = csr_mstatus_mie;
            csr_mstatus_mie_nxt = 0;
            csr_mstatus_mpp_nxt = csr_mcurrent_privilege;
            csr_mcurrent_privilege_nxt = `ARMLEOCPU_PRIVILEGE_MACHINE;

            csr_mepc_nxt = csr_exc_epc;
            csr_next_pc = csr_mtvec;
        end
    end else if((csr_cmd == `ARMLEOCPU_CSR_CMD_MRET) && (csr_mcurrent_privilege_machine)) begin
        csr_mstatus_mie_nxt = csr_mstatus_mpie;
        csr_mstatus_mpie_nxt = 1;
        csr_mstatus_mprv_nxt = 0; // Changed in v1.12 of privileged spec

        csr_next_pc = csr_mepc;
        csr_cmd_exc_int_error = 0;
    end else if(csr_cmd == `ARMLEOCPU_CSR_CMD_SRET && (csr_mcurrent_privilege_machine_supervisor)) begin
        csr_mstatus_sie_nxt = csr_mstatus_spie;
        csr_mstatus_spie_nxt = 1;
        csr_mstatus_mprv_nxt = 0; // Changed in v1.12 of privileged spec

        csr_next_pc = csr_sepc;
        csr_cmd_exc_int_error = 0;
    end else if(csr_cmd == `ARMLEOCPU_CSR_CMD_EXCEPTION_BEGIN) begin
        csr_mstatus_mpie_nxt = csr_mstatus_mie;
        csr_mstatus_mie_nxt = 0;
        csr_mstatus_mpp_nxt = csr_mcurrent_privilege;
        csr_mcurrent_privilege_nxt = `ARMLEOCPU_PRIVILEGE_MACHINE;
        csr_mepc_nxt = csr_exc_epc;
        csr_next_pc = csr_mtvec;
        

        csr_mcause_nxt = csr_exc_cause;
        csr_cmd_exc_int_error = 0;
    end else if(csr_write || csr_read) begin
        csr_cmd_exc_int_error = 0;
        case(csr_address)
            `DEFINE_CSR_COMB_RO(12'hF11, MVENDORID)
            `DEFINE_CSR_COMB_RO(12'hF12, MARCHID)
            `DEFINE_CSR_COMB_RO(12'hF13, MIMPID)
            `DEFINE_CSR_COMB_RO(12'hF14, MHARTID)
            // Added in v1.12
            `DEFINE_CSR_COMB_RO(12'hF15, MCONFIGPTR)
            12'hBC0: begin // MCURRENT_PRIVILEGE
                // This is used only for debug purposes
                // TODO: Fix this to bne readonly
                csr_exists = 1;
                csr_to_rd = {30'h0, csr_mcurrent_privilege};
                rmw_before = csr_to_rd;
                if(!csr_invalid && csr_write && (rmw_after[1:0] != 2'b10)) begin
                    csr_mcurrent_privilege_nxt = rmw_after[1:0];
                end
            end
            12'h300: begin // MSTATUS
                csr_exists = 1;
                csr_to_rd = {
                            9'h0, // Padding SD, 8 empty bits
                            csr_mstatus_tsr, csr_mstatus_tw, csr_mstatus_tvm, // trap enable bits
                            csr_mstatus_mxr, csr_mstatus_sum, csr_mstatus_mprv, //machine privilege mode
                            2'b00, 2'b00, // xs, fs
                            csr_mstatus_mpp, 2'b00, csr_mstatus_spp, // MPP, 2 bits (reserved by spec), SPP
                            csr_mstatus_mpie, 1'b0, csr_mstatus_spie, 1'b0,
                            csr_mstatus_mie, 1'b0, csr_mstatus_sie, 1'b0};
                rmw_before = csr_to_rd;
                if(!csr_invalid && csr_write) begin
                    csr_mstatus_tsr_nxt = rmw_after[22];
                    csr_mstatus_tw_nxt = rmw_after[21];
                    csr_mstatus_tvm_nxt = rmw_after[20];
                    csr_mstatus_mxr_nxt = rmw_after[19];
                    csr_mstatus_sum_nxt = rmw_after[18];
                    csr_mstatus_mprv_nxt = rmw_after[17];

                    if(rmw_after[12:11] != 2'b10)
                        csr_mstatus_mpp_nxt = rmw_after[12:11];
                    csr_mstatus_spp_nxt = rmw_after[8];

                    csr_mstatus_mpie_nxt = rmw_after[7];
                    csr_mstatus_spie_nxt = rmw_after[5];
                    csr_mstatus_mie_nxt = rmw_after[3];
                    csr_mstatus_sie_nxt = rmw_after[1];
                end
            end
            // MSTATUSH
            // Added in v1.12 of privileged spec
            `DEFINE_CSR_COMB_RO(12'h310, 0)

            `DEFINE_CSR_COMB_RO(12'h301, csr_misa)

            //Intentionally not implemented: `DEFINE_CSR_COMB_RO(12'h320, 0) // mcountinhibit

            `DEFINE_CSR_COMB_RO(12'h306, 0) // mcounteren

            `DEFINE_CSR_COMB_RO(12'h106, 0) // scounteren


            // Value should be written for all valid bits, and invalids are ignored
            // Also note that *TVEC CSR may change in future
            // Because 2 bottom bits are used to select interrupt scheme

            `DEFINE_ADDRESS_CSR_REG_COMB(12'h305, csr_mtvec)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'h340, csr_mscratch)
            `DEFINE_ADDRESS_CSR_REG_COMB(12'h341, csr_mepc)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'h342, csr_mcause)
            `DEFINE_CSR_COMB_RO(12'h343, 0)
            // MTVAL is hardwired to zero, in case it never gets written
            
            // Supervisor
            `DEFINE_ADDRESS_CSR_REG_COMB(12'h105, csr_stvec)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'h140, csr_sscratch)
            `DEFINE_ADDRESS_CSR_REG_COMB(12'h141, csr_sepc)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'h142, csr_scause)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'h143, csr_stval)
            // STVAL is NOT hardwired to zero
            

            `DEFINE_SCRATCH_CSR_REG_COMB(12'hB00, csr_cycle)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'hB80, csr_cycleh)

            `DEFINE_SCRATCH_CSR_REG_COMB(12'hB02, csr_instret)
            `DEFINE_SCRATCH_CSR_REG_COMB(12'hB82, csr_instreth)
            12'h180: begin // SATP
                csr_to_rd = {csr_satp_mode, 9'h0, csr_satp_ppn};
                csr_exists = !(csr_mstatus_tvm && csr_mcurrent_privilege_supervisor);
                rmw_before = csr_to_rd;
                if(!csr_invalid && csr_write) begin
                    csr_satp_mode_nxt = rmw_after[31];
                    csr_satp_ppn_nxt = rmw_after[21:0];
                end
            end
            // MEDELEG
            `DEFINE_CSR_COMB_RO(12'h302, 0)
            // MIDELEG
            `DEFINE_CSR_COMB_RO(12'h303, 0)

            12'h304: begin // MIE
                csr_exists = 1;

                csr_to_rd[11] = csr_mie_meie;
                csr_to_rd [9] = csr_mie_seie;

                csr_to_rd [7] = csr_mie_mtie;
                csr_to_rd [5] = csr_mie_stie;

                csr_to_rd [3] = csr_mie_msie;
                csr_to_rd [1] = csr_mie_ssie;

                rmw_before = csr_to_rd;
                if(csr_write && !csr_invalid) begin
                    csr_mie_meie_nxt = rmw_after[11];
                    csr_mie_seie_nxt = rmw_after [9];
                    csr_mie_mtie_nxt = rmw_after [7];
                    csr_mie_stie_nxt = rmw_after [5];
                    csr_mie_msie_nxt = rmw_after [3];
                    csr_mie_ssie_nxt = rmw_after [1];
                end
            end
            12'h104: begin // SIE
                csr_exists = 1;
                csr_to_rd [9] = csr_mie_seie;

                csr_to_rd [5] = csr_mie_stie;

                csr_to_rd [1] = csr_mie_ssie;

                rmw_before = csr_to_rd;
                if(!csr_invalid && csr_write) begin
                    csr_mie_seie_nxt = rmw_after [9];
                    csr_mie_stie_nxt = rmw_after [5];
                    csr_mie_ssie_nxt = rmw_after [1];
                end
            end
            12'h100: begin // SSTATUS
                csr_exists = 1;
                csr_to_rd = {
                            9'h0, // Padding SD, 9 empty bits
                            3'b000, // trap enable bits
                            csr_mstatus_mxr, csr_mstatus_sum, 1'b0, //mxr, sum, mprv
                            2'b00, 2'b00, // xs, fs
                            2'b00, 2'b00, csr_mstatus_spp, // MPP, 2 bits (reserved by spec), SPP
                            1'b0, 1'b0, csr_mstatus_spie, 1'b0,
                            1'b0, 1'b0, csr_mstatus_sie, 1'b0};
                rmw_before = csr_to_rd;
                if(!csr_invalid && csr_write) begin
                    csr_mstatus_mxr_nxt = rmw_after[19];
                    csr_mstatus_sum_nxt = rmw_after[18];
                    csr_mstatus_spp_nxt = rmw_after[8];
                    csr_mstatus_spie_nxt = rmw_after[5];
                    csr_mstatus_sie_nxt = rmw_after[1];
                end
            end
            
            12'h344: begin // MIP
                csr_exists = 1;
                rmw_before = 0;

                // meip
                // 11th bit, read only
                rmw_before[11] = irq_meip_i;

                // s*ip bit, read/write
                // when read s*ip is logical or of this bit and external signal
                // when rmw then s*ip is this bit
                
                rmw_before[9] = csr_mip_seip;
                

                // TIMER
                rmw_before[7] = irq_mtip_i;
                
                rmw_before[5] = csr_mip_stip;
                
                // SWI
                rmw_before[3] = irq_msip_i;
                
                rmw_before[1] = csr_mip_ssip;

                // We write to rd the value ored with external input
                // But we only RMW the saved register value
                csr_to_rd = rmw_before;

                // s*ip bit, read/write
                // when read seip is logical or of this bit and external signal
                // when rmw then seip is this bit
            
                csr_to_rd[9] = irq_calculated_seip;
                
                csr_to_rd[5] = irq_calculated_stip;
                
                csr_to_rd[1] = irq_calculated_ssip;
                

                if(!csr_invalid && csr_write) begin
                    // csr_mip_m*ip is read only

                    csr_mip_seip_nxt = rmw_after[9];
                
                    csr_mip_stip_nxt = rmw_after[5];
                
                    csr_mip_ssip_nxt = rmw_after[1];
                end
            end
            12'h144: begin // SIP
                csr_exists = 1;

                // s*ip bit, read/write
                // when read seip is logical or of this bit and external signal
                // when rmw then seip is this bit
                
                rmw_before[9] = csr_mip_seip;
                
                rmw_before[5] = csr_mip_stip;
                
                rmw_before[1] = csr_mip_ssip;


                csr_to_rd = rmw_before;

                csr_to_rd[9] = irq_calculated_seip;
                
                csr_to_rd[5] = irq_calculated_stip;
                
                csr_to_rd[1] = irq_calculated_ssip;
                
                if(!csr_invalid && csr_write) begin
                    // csr_mip_m*ip is read only
                    csr_mip_seip_nxt = rmw_after[9];
                    
                    csr_mip_stip_nxt = rmw_after[5];
                    
                    csr_mip_ssip_nxt = rmw_after[1];
                end
            end
            
            default: begin
                // By default in logic above
                // csr_exists = 0;
                // and all rmw and csr_to_rd is set to zero

                // For HPM COUNTER
                if((csr_address >= 12'hB03) && (csr_address <= 12'hB1F)) begin
                    csr_exists = 1;
                    // Pretend it exists and is hardwired to zero
                end
                // For HPM COUNTER High section
                if((csr_address >= 12'hB83) && (csr_address <= 12'hB9F)) begin
                    csr_exists = 1;
                    // Pretend it exists and is hardwired to zero
                end
                // For HPM EVENT registers
                if((csr_address >= 12'h323) && (csr_address <= 12'h33F)) begin
                    csr_exists = 1;
                    // Pretend it exists and is hardwired to zero
                end
                
                
            end
        endcase
    end else if(csr_cmd == `ARMLEOCPU_CSR_CMD_NONE) begin
        csr_cmd_exc_int_error = 0;
    end // else csr_cmd_exc_int_error = 1; but no need because it's 1 by default
end



`ifdef FORMAL_RULES
// verilator coverage_off
    always @(posedge clk) begin
        if(csr_cmd == `ARMLEOCPU_CSR_CMD_MRET)
            assert(csr_mcurrent_privilege_machine);
        if(csr_cmd == `ARMLEOCPU_CSR_CMD_SRET)
            assert(
                (csr_mcurrent_privilege_machine)
                || (csr_mcurrent_privilege_supervisor));
    end
// verilator coverage_on
`endif

// TODO: Add logging

endmodule

`include "armleocpu_undef.vh"
