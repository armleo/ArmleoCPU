// ALU_OUTPUT_SELECT
`define ALU_SELECT_ADD 4'd0
`define ALU_SELECT_SUB 4'd1
`define ALU_SELECT_SLT 4'd2
`define ALU_SELECT_SLTU 4'd3
`define ALU_SELECT_SLL 4'd4
`define ALU_SELECT_SRA 4'd5
`define ALU_SELECT_SRL 4'd6
`define ALU_SELECT_XOR 4'd7
`define ALU_SELECT_OR 4'd8
`define ALU_SELECT_AND 4'd9

`define ALU_SELECT_WIDTH 4

// ARMLEOBUS
`define ARMLEOBUS_CMD_NONE (3'd0)
`define ARMLEOBUS_CMD_READ (3'd1)
`define ARMLEOBUS_CMD_WRITE (3'd2)

`define ARMLEOBUS_RESPONSE_SUCCESS (3'd0)
`define ARMLEOBUS_UNKNOWN_ADDRESS (3'd1)
`define ARMLEOBUS_INVALID_OPERATION (3'd2)

// ACCESSTAG
`define ACCESSTAG_W (8)

`define ACCESSTAG_VALID_BIT_NUM (0)
`define ACCESSTAG_READ_BIT_NUM (1)
`define ACCESSTAG_WRITE_BIT_NUM (2)
`define ACCESSTAG_EXECUTE_BIT_NUM (3)
`define ACCESSTAG_USER_BIT_NUM (4)
`define ACCESSTAG_ACCESS_BIT_NUM (6)
`define ACCESSTAG_DIRTY_BIT_NUM (7)

// CACHE
`define CACHE_RESPONSE_IDLE (4'd0)
`define CACHE_RESPONSE_WAIT (4'd1)
`define CACHE_RESPONSE_DONE (4'd2)
`define CACHE_RESPONSE_ACCESSFAULT (4'd3)
`define CACHE_RESPONSE_PAGEFAULT (4'd4)
`define CACHE_RESPONSE_MISSALIGNED (4'd5)
`define CACHE_RESPONSE_UNKNOWNTYPE (4'd6)

`define CACHE_CMD_NONE (4'd0)
`define CACHE_CMD_EXECUTE (4'd1)
`define CACHE_CMD_LOAD (4'd2)
`define CACHE_CMD_STORE (4'd3)
`define CACHE_CMD_FLUSH_ALL (4'd4)

`define CACHE_ERROR_ACCESSFAULT (1'd0)
`define CACHE_ERROR_PAGEFAULT (1'd1)

// CSR CMDs

`define ARMLEOCPU_CSR_CMD_NONE (4'd0)
`define ARMLEOCPU_CSR_CMD_READ (4'd1)
`define ARMLEOCPU_CSR_CMD_WRITE (4'd2)
`define ARMLEOCPU_CSR_CMD_READ_WRITE (4'd3)
`define ARMLEOCPU_CSR_CMD_READ_SET (4'd4)
`define ARMLEOCPU_CSR_CMD_READ_CLEAR (4'd5)
`define ARMLEOCPU_CSR_CMD_MRET (4'd6)
`define ARMLEOCPU_CSR_CMD_SRET (4'd7)
`define ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN (4'd8)

// E2F CMDs
`define ARMLEOCPU_E2F_CMD_WIDTH 3
`define ARMLEOCPU_E2F_CMD_BUBBLE_JUMP (3'h3)
`define ARMLEOCPU_E2F_CMD_FLUSH (3'h2)
`define ARMLEOCPU_E2F_CMD_BRANCHTAKEN (3'h1)
`define ARMLEOCPU_E2F_CMD_IDLE (3'h0)


// Exceptions and interrupts
`define EXCEPTION_CODE_INTERRUPT (32'h8000_0000)
`define INTERRUPT_CODE_SOFTWATE_INTERRUPT (3)
`define INTERRUPT_CODE_TIMER_INTERRUPT (7)
`define INTERRUPT_CODE_EXTERNAL_INTERRUPT (11)

`define EXCEPTION_CODE_SOFTWATE_INTERRUPT (`INTERRUPT_CODE_SOFTWATE_INTERRUPT | `EXCEPTION_CODE_INTERRUPT)
`define EXCEPTION_CODE_TIMER_INTERRUPT (`INTERRUPT_CODE_TIMER_INTERRUPT | `EXCEPTION_CODE_INTERRUPT)
`define EXCEPTION_CODE_EXTERNAL_INTERRUPT (`INTERRUPT_CODE_EXTERNAL_INTERRUPT | `EXCEPTION_CODE_INTERRUPT)

`define EXCEPTION_CODE_INSTRUCTION_ADDRESS_MISSALIGNED (0)
`define EXCEPTION_CODE_INSTRUCTION_ACCESS_FAULT (1)
`define EXCEPTION_CODE_ILLEGAL_INSTRUCTION (2)
`define EXCEPTION_CODE_BREAKPOINT (3)
`define EXCEPTION_CODE_LOAD_ADDRESS_MISALIGNED (4)
`define EXCEPTION_CODE_LOAD_ACCESS_FAULT (5)
`define EXCEPTION_CODE_STORE_ADDRESS_MISALIGNED (6)
`define EXCEPTION_CODE_STORE_ACCESS_FAULT (7)

// Calls from x privilege
`define EXCEPTION_CODE_UCALL (8)
`define EXCEPTION_CODE_SCALL (9)
`define EXCEPTION_CODE_MCALL (11)
`define EXCEPTION_CODE_INSTRUCTION_PAGE_FAULT (12)
`define EXCEPTION_CODE_LOAD_PAGE_FAULT (13)
`define EXCEPTION_CODE_STORE_PAGE_FAULT (15)


// INSTRs
`define INSTRUCTION_NOP ({12'h0, 5'h0, 3'b000, 5'h0, 7'b00_100_11})

`define OPCODE_LUI (7'b0110111)
`define OPCODE_AUIPC (7'b0010111)
`define OPCODE_JAL (7'b1101111)
`define OPCODE_JALR (7'b1100111)
`define OPCODE_BRANCH (7'b1100011)
`define OPCODE_LOAD (7'b0000011)
`define OPCODE_STORE (7'b0100011)
`define OPCODE_OP_IMM (7'b0010011)
`define OPCODE_OP (7'b0110011)
`define OPCODE_FENCE (7'b0001111)
`define OPCODE_SYSTEM (7'b1110011)

// Privileges
`define ARMLEOCPU_PRIVILEGE_USER (2'b00)
`define ARMLEOCPU_PRIVILEGE_USER_SV (1'b0)
`define ARMLEOCPU_PRIVILEGE_SUPERVISOR (2'b01)
`define ARMLEOCPU_PRIVILEGE_SUPERVISOR_SV (1'b1)
`define ARMLEOCPU_PRIVILEGE_MACHINE (2'b11)

// TLB CMDs
`define TLB_CMD_NONE (2'b00)
`define TLB_CMD_RESOLVE (2'b01)
`define TLB_CMD_WRITE (2'b10)
`define TLB_CMD_INVALIDATE (2'b11)


// LD_TYOE
`define LOAD_BYTE (3'b000)
`define LOAD_BYTE_UNSIGNED (3'b100)

`define LOAD_HALF (3'b001)
`define LOAD_HALF_UNSIGNED (3'b101)

`define LOAD_WORD (3'b010)

// ST_TYPE
`define STORE_BYTE (2'b00)
`define STORE_HALF (2'b01)
`define STORE_WORD (2'b10)
