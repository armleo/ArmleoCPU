module armleocpu_control(
    
);

endmodule