
localparam ACCESSTAG_W = 8;

localparam OPCODE_LUI    = 7'b0110111;
localparam OPCODE_AUIPC  = 7'b0010111;
localparam OPCODE_JAL    = 7'b1101111;
localparam OPCODE_JALR   = 7'b1100111;
localparam OPCODE_BRANCH = 7'b1100011;
localparam OPCODE_LOAD   = 7'b0000011;
localparam OPCODE_STORE  = 7'b0100011;
localparam OPCODE_ALUI   = 7'b0010011;
localparam OPCODE_ALU    = 7'b0110011;
localparam OPCODE_MISCMEM= 7'b0001111;
localparam OPCODE_SYSTEM = 7'b1110011;


localparam EXCEPTION_CODE_INTERRUPT = 32'h8000_0000;
localparam EXCEPTION_CODE_SOFTWATE_INTERRUPT = 3 | EXCEPTION_CODE_INTERRUPT;
localparam EXCEPTION_CODE_TIMER_INTERRUPT = 7 | EXCEPTION_CODE_INTERRUPT;
localparam EXCEPTION_CODE_EXTERNAL_INTERRUPT = 11 | EXCEPTION_CODE_INTERRUPT;

localparam EXCEPTION_CODE_INSTRUCTION_ADDRESS_MISALIGNED = 0;
localparam EXCEPTION_CODE_INSTRUCTION_ACCESS_FAULT = 1;
localparam EXCEPTION_CODE_ILLEGAL_INSTRUCTION = 2;
localparam EXCEPTION_CODE_BREAKPOINT = 3;
localparam EXCEPTION_CODE_LOAD_ADDRESS_MISALIGNED = 4;
localparam EXCEPTION_CODE_LOAD_ACCESS_FAULT = 5;
localparam EXCEPTION_CODE_STORE_ADDRESS_MISALIGNED = 6;
localparam EXCEPTION_CODE_STORE_ACCESS_FAULT = 7;

// Calls from x privilege
localparam EXCEPTION_CODE_UCALL = 8;
localparam EXCEPTION_CODE_SCALL = 9;
localparam EXCEPTION_CODE_MCALL = 11;
localparam EXCEPTION_CODE_INSTRUCTION_PAGE_FAULT = 12;
localparam EXCEPTION_CODE_LOAD_PAGE_FAULT = 13;
localparam EXCEPTION_CODE_STORE_PAGE_FAULT = 15;



// ST_TYPE
localparam STORE_BYTE = 2'b00;
localparam STORE_HALF = 2'b01;
localparam STORE_WORD = 2'b10;


// LD_TYPE
localparam LOAD_BYTE = 3'b000;
localparam LOAD_BYTE_UNSIGNED = 3'b100;

localparam LOAD_HALF = 3'b001;
localparam LOAD_HALF_UNSIGNED = 3'b101;

localparam LOAD_WORD = 3'b010;


localparam CACHE_RESPONSE_WAIT        = 3'd0;
localparam CACHE_RESPONSE_DONE        = 3'd1;
localparam CACHE_RESPONSE_ACCESSFAULT = 3'd2;
localparam CACHE_RESPONSE_PAGEFAULT   = 3'd3;
localparam CACHE_RESPONSE_MISSALIGNED = 3'd4;
localparam CACHE_RESPONSE_UNKNOWNTYPE = 3'd5;

localparam ACCESSTAG_VALID_BIT_NUM = 0;
localparam ACCESSTAG_READ_BIT_NUM = 1;
localparam ACCESSTAG_WRITE_BIT_NUM = 2;
localparam ACCESSTAG_EXECUTE_BIT_NUM = 3;
localparam ACCESSTAG_USER_BIT_NUM = 4;
localparam ACCESSTAG_ACCESS_BIT_NUM = 6;
localparam ACCESSTAG_DIRTY_BIT_NUM = 7;





