
// ST_TYPE
localparam STORE_BYTE = 2'b00;
localparam STORE_HALF = 2'b01;
localparam STORE_WORD = 2'b10;
