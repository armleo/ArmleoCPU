`define CACHE_RESPONSE_WAIT 3'd0
`define CACHE_RESPONSE_DONE 3'd1
`define CACHE_RESPONSE_ACCESSFAULT 3'd2
`define CACHE_RESPONSE_PAGEFAULT 3'd3
`define CACHE_RESPONSE_MISSALIGNED 3'd4
`define CACHE_RESPONSE_UNKNOWNTYPE 3'd5

`define CACHE_CMD_NONE 3'd0
`define CACHE_CMD_EXECUTE 3'd1
`define CACHE_CMD_LOAD 3'd2
`define CACHE_CMD_STORE 3'd3
`define CACHE_CMD_FLUSH 3'd4


