
`define ACCESSTAG_W (8)

`define ACCESSTAG_VALID_BIT_NUM (0)
`define ACCESSTAG_READ_BIT_NUM (1)
`define ACCESSTAG_WRITE_BIT_NUM (2)
`define ACCESSTAG_EXECUTE_BIT_NUM (3)
`define ACCESSTAG_USER_BIT_NUM (4)
`define ACCESSTAG_ACCESS_BIT_NUM (6)
`define ACCESSTAG_DIRTY_BIT_NUM (7)





