`define DECODE_IS_OP_IMM 0
`define DECODE_IS_OP 1
`define DECODE_IS_JALR 2
`define DECODE_IS_JAL 3
`define DECODE_IS_LUI 4
`define DECODE_IS_AUIPC 5
`define DECODE_IS_BRANCH 6
`define DECODE_IS_STORE 7
`define DECODE_IS_LOAD 8


`define DECODE_IS_MUL 9
`define DECODE_IS_MULH 10
`define DECODE_IS_MULHSU 11
`define DECODE_IS_MULHU 12

`define DECODE_IS_DIV 13
`define DECODE_IS_DIVU 14

`define DECODE_IS_REM 15
`define DECODE_IS_REMU 16

`define DECODE_IS_EBREAK 17

`define DECODE_IS_ECALL 18
`define DECODE_IS_WFI 19
`define DECODE_IS_MRET 20
`define DECODE_IS_SRET 21

`define DECODE_IS_SFENCE_VMA 22
`define DECODE_IS_IFENCEI 23

`define DECODE_IS_FENCE_NORMAL 24

`define DECODE_IS_CSRRW_CSRRWI 25
`define DECODE_IS_CSRS_CSRSI 26
`define DECODE_IS_CSRC_CSRCI 27

`define DECODE_IS_CSR 28

// contains decode's output length
`define DECODE_IS_WIDTH 29



`define OPCODE_LUI (7'b0110111)
`define OPCODE_AUIPC (7'b0010111)
`define OPCODE_JAL (7'b1101111)
`define OPCODE_JALR (7'b1100111)
`define OPCODE_BRANCH (7'b1100011)
`define OPCODE_LOAD (7'b0000011)
`define OPCODE_STORE (7'b0100011)
`define OPCODE_OP_IMM (7'b0010011)
`define OPCODE_OP (7'b0110011)
`define OPCODE_FENCE (7'b0001111)
`define OPCODE_SYSTEM (7'b1110011)