
localparam ACCESSTAG_W = 8;

localparam ACCESSTAG_VALID_BIT_NUM = 0;
localparam ACCESSTAG_READ_BIT_NUM = 1;
localparam ACCESSTAG_WRITE_BIT_NUM = 2;
localparam ACCESSTAG_EXECUTE_BIT_NUM = 3;
localparam ACCESSTAG_USER_BIT_NUM = 4;
localparam ACCESSTAG_ACCESS_BIT_NUM = 6;
localparam ACCESSTAG_DIRTY_BIT_NUM = 7;





