
`define ARMLEOBUS_CMD_NONE 3'd0
`define ARMLEOBUS_CMD_READ 3'd1
`define ARMLEOBUS_CMD_WRITE 3'd2

`define ARMLEOBUS_RESPONSE_SUCCESS 3'd0
`define ARMLEOBUS_UNKNOWN_ADDRESS 3'd1
`define ARMLEOBUS_INVALID_OPERATION 3'd2

