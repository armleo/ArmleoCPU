

// LD_TYPE
localparam LOAD_BYTE = 3'b000;
localparam LOAD_BYTE_UNSIGNED = 3'b100;

localparam LOAD_HALF = 3'b001;
localparam LOAD_HALF_UNSIGNED = 3'b101;

localparam LOAD_WORD = 3'b010;
