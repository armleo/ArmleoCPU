module armleocpu_execute(
    input clk,
    input rst_n,

// Fetch unit
    input      [31:0]       f2e_instr,
    input      [31:0]       f2e_pc,
    input                   f2e_exc_start,
    input                   f2e_exc_return,
    input      [1:0]        f2e_exc_privilege,
    input      [31:0]       f2e_epc,
    input      [31:0]       f2e_cause,

    output reg              e2f_ready,
    output reg  [1:0]       e2f_cmd,
    output reg [31:0]       e2f_bubble_exc_start_target,
    output reg [31:0]       e2f_bubble_exc_return_target,
    output reg [31:0]       e2f_branchtarget,

// To debug unit, indicates that ebreak in machine mode was met
    output reg              e2debug_machine_ebreak,

// Cache interface
    input      [3:0]        c_response,
    input                   c_reset_done,

    output reg [3:0]        c_cmd,
    output reg [31:0]       c_address,
    output     [2:0]        c_load_type,
    input      [31:0]       c_load_data,
    output     [1:0]        c_store_type,
    output     [31:0]       c_store_data,


// CSR Interface for csr class instructions
    output reg [3:0]        csr_cmd, // NONE, WRITE, READ, READ_WRITE, 
    output     [11:0]       csr_address,
    input                   csr_invalid,
    input      [31:0]       csr_readdata,
    output reg [31:0]       csr_writedata,

    input      [31:0]       csr_next_pc,
    output     [31:0]       csr_exc_cause,
    output     [31:0]       csr_exc_epc,
    output     [1:0]        csr_exc_privilege,

// CSR Registers
    input      [1:0]        csr_mcurrent_privilege,
    input      [31:0]       csr_mepc,
    input      [31:0]       csr_sepc,
    
    input                   csr_mstatus_tsr, // sret generates illegal instruction
    input                   csr_mstatus_tvm, // sfence vma and csr satp write generates illegal instruction
    input                   csr_mstatus_tw, // wfi generates illegal instruction

// Regfile
    output     [4:0]        rs1_addr,
    input      [31:0]       rs1_data,

    output     [4:0]        rs2_addr,
    input      [31:0]       rs2_data,
    
    output     [4:0]        rd_addr,
    output reg [31:0]       rd_wdata,
    output reg              rd_write
);

`include "armleocpu_cache.vh"
`include "armleocpu_instructions.vh"
`include "armleocpu_exception.vh"
`include "armleocpu_privilege.vh"
`include "armleocpu_csr.vh"

// |------------------------------------------------|
// |              State                             |
// |------------------------------------------------|

reg dcache_command_issued;
reg csr_done;

// |------------------------------------------------|
// |              Signals                           |
// |------------------------------------------------|

// Decode opcode
wire [6:0]  opcode                  = f2e_instr[6:0];
assign      rd_addr                 = f2e_instr[11:7];
wire [2:0]  funct3                  = f2e_instr[14:12];
assign      rs1_addr                = f2e_instr[19:15];
assign      rs2_addr                = f2e_instr[24:20];
wire [6:0]  funct7                  = f2e_instr[31:25];
assign      c_load_type             = funct3;
assign      c_store_type            = funct3[1:0];
assign      c_store_data            = rs2_data;

//
//
//
wire sign = f2e_instr[31];

wire [31:0] immgen_simm12 = {{20{sign}}, f2e_instr[31:20]};
wire [31:0] immgen_store_offset = {{20{sign}}, f2e_instr[31:25], f2e_instr[11:7]};
wire [31:0] immgen_branch_offset = {{20{sign}}, f2e_instr[7], f2e_instr[30:25], f2e_instr[11:8], 1'b0};
wire [31:0] immgen_upper_imm = {f2e_instr[31:12], 12'h000};
wire [31:0] immgen_jal_offset = {{12{sign}}, f2e_instr[19:12], f2e_instr[20], f2e_instr[30:25], f2e_instr[24:21], 1'b0};
// 11 + 1 + 6 + 1 + 6 + 4 + 1
wire [31:0] immgen_csr_imm = {27'b0, f2e_instr[19:15]}; // used by csr bit write/set/clear


assign      csr_exc_epc             = f2e_pc;

wire is_op_imm  = opcode == `OPCODE_OP_IMM;
wire is_op      = opcode == `OPCODE_OP;
wire is_jalr    = opcode == `OPCODE_JALR;
wire is_jal     = opcode == `OPCODE_JAL;
wire is_lui     = opcode == `OPCODE_LUI;
wire is_auipc   = opcode == `OPCODE_AUIPC;
wire is_branch  = opcode == `OPCODE_BRANCH;
wire is_store   = opcode == `OPCODE_STORE;
wire is_load    = opcode == `OPCODE_LOAD;
wire is_system  = opcode == `OPCODE_SYSTEM;
wire is_fence   = opcode == `OPCODE_FENCE;

wire is_ebreak  = f2e_instr == 32'b000000000001_00000_000_00000_1110011;

wire is_mul         = is_op     && (funct3 == 3'b000) && (funct7 == 7'b0000_001);
wire is_mulh        = is_op     && (funct3 == 3'b001) && (funct7 == 7'b0000_001);
wire is_mulhsu      = is_op     && (funct3 == 3'b010) && (funct7 == 7'b0000_001);
wire is_mulhu       = is_op     && (funct3 == 3'b011) && (funct7 == 7'b0000_001);

wire is_div         = is_op     && (funct3 == 3'b100) && (funct7 == 7'b0000_001);
wire is_divu        = is_op     && (funct3 == 3'b101) && (funct7 == 7'b0000_001);

wire is_rem         = is_op     && (funct3 == 3'b110) && (funct7 == 7'b0000_001);
wire is_remu        = is_op     && (funct3 == 3'b111) && (funct7 == 7'b0000_001);


wire dcache_response_done = c_response == `CACHE_RESPONSE_DONE;
wire dcache_response_error = (c_response == `CACHE_RESPONSE_MISSALIGNED) || (c_response == `CACHE_RESPONSE_ACCESSFAULT) || (c_response == `CACHE_RESPONSE_PAGEFAULT);
// TODO:

reg illegal_instruction;
reg dcache_exc;
reg [31:0] dcache_exc_cause;


wire [31:0] alu_result;
wire alu_illegal_instruction;

wire [31:0] pc_plus_4 = f2e_pc + 4;

wire brcond_branchtaken;
wire brcond_illegal_instruction;

reg mul_valid;
reg [31:0] mul_factor0;
reg [31:0] mul_factor1;

wire mul_ready;
wire [63:0] mul_result;
wire [63:0] mul_inverted_result = -mul_result;

reg div_fetch;
reg div_signinvert;
reg [31:0] div_dividend;
reg [31:0] div_divisor;

wire div_ready;
wire div_division_by_zero;
wire [31:0] div_quotient;
wire [31:0] div_remainder;

// |------------------------------------------------|
// |              ALU                               |
// |------------------------------------------------|
armleocpu_alu alu(
    .is_op_imm(is_op_imm),
    .is_op(is_op),

    .funct3(funct3),
    .funct7(funct7),
    .shamt(f2e_instr[24:20]),

    .rs1(rs1_data),
    .rs2(rs2_data),
    
    .simm12(immgen_simm12),

    .result(alu_result),
    .illegal_instruction(alu_illegal_instruction)
);

// |------------------------------------------------|
// |              brcond                               |
// |------------------------------------------------|
armleocpu_brcond brcond(
    .funct3                 (funct3),
    .rs1                    (rs1_data),
    .rs2                    (rs2_data),
    .incorrect_instruction  (brcond_illegal_instruction),
    .branch_taken           (brcond_branchtaken)
);

armleocpu_multiplier multiplier(
    .clk            (clk),
    .rst_n          (rst_n),

    .valid          (mul_valid),

    .factor0        (mul_factor0),
    .factor1        (mul_factor1),

    .ready          (mul_ready),
    .result         (mul_result)
);


armleocpu_unsigned_divider divider(
    .clk                (clk),
    .rst_n              (rst_n),

    .fetch              (div_fetch),

    .dividend           (div_dividend),
    .divisor            (div_divisor),

    .ready              (div_ready),
    .division_by_zero   (div_division_by_zero),
    .quotient           (div_quotient),
    .remainder          (div_remainder)        
);
reg [3:0] rd_sel;
reg mul_signinvert;
`define RD_ALU (4'd0)
`define RD_CSR (4'd1)
`define RD_DCACHE (4'd2)
`define RD_LUI (4'd3)
`define RD_AUIPC (4'd4)
`define RD_PC_PLUS_4 (4'd5)
`define RD_MUL (4'd6)
`define RD_MULH (4'd7)
`define RD_DIV (4'd8)
`define RD_REM (4'd9)
`define RD_RS1 (4'd10)
`define RD_MINUS_ONE (4'd11)

always @* begin
    case(rd_sel)
        `RD_ALU:        rd_wdata = alu_result;
        `RD_CSR:        rd_wdata = csr_readdata;
        `RD_DCACHE:     rd_wdata = c_load_data;
        `RD_LUI:        rd_wdata = immgen_upper_imm;
        `RD_AUIPC:      rd_wdata = f2e_pc + immgen_upper_imm;
        `RD_PC_PLUS_4:  rd_wdata = pc_plus_4;
        `RD_MUL:        rd_wdata = mul_signinvert ? mul_inverted_result[31:0] : mul_result[31:0];
        `RD_MULH:       rd_wdata = mul_signinvert ? mul_inverted_result[63:32] : mul_result[63:32];
        `RD_DIV:        rd_wdata = div_signinvert ? -div_quotient : div_quotient;
        `RD_REM:        rd_wdata = div_signinvert ? -div_remainder : div_remainder;
        `RD_RS1:        rd_wdata = rs1_data;
        `RD_MINUS_ONE:  rd_wdata = -1;
        default:        rd_wdata = alu_result;
    endcase
end

// TODO:
// assign e2f_bubble_exc_start_target = ;

always @* begin
    illegal_instruction = 0;
    e2f_ready = 1;
    e2f_branchtarget = f2e_pc + immgen_branch_offset;
    e2f_cmd = `ARMLEOCPU_E2F_CMD_IDLE;
    e2f_bubble_exc_start_target = csr_next_pc;
    e2f_bubble_exc_return_target = csr_next_pc;

    e2debug_machine_ebreak = 0;

    c_cmd = `CACHE_CMD_NONE;
    c_address = rs1_data + immgen_simm12;
    

    csr_cmd = `CSR_CMD_NONE;
    csr_writedata = 0;
    csr_exc_cause = 20;
    csr_exc_epc = csr_mepc;
    csr_exc_privilege = `ARMLEOCPU_PRIVILEGE_USER;

    rd_write = 0;
    mul_signinvert = 0;

    rd_sel = `RD_ALU;
    
    dcache_exc = 0;
    dcache_exc_cause = 0;

    mul_valid = 0;

    mul_factor0 = rs1_data;
    mul_factor1 = rs2_data;

    div_fetch = 0;
    div_signinvert = 0;
    div_dividend = rs1_data;
    div_divisor = rs2_data;

    case(1)
        is_mul: begin
            e2f_ready = 0;
            mul_signinvert = rs1_data[31] ^ rs2_data[31];
            mul_valid = !mul_ready;
            mul_factor0 = rs1_data[31] ? -rs1_data : rs1_data;
            mul_factor1 = rs2_data[31] ? -rs2_data : rs2_data;
            if(mul_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_MUL;
            end
        end
        is_mulh: begin
            e2f_ready = 0;
            mul_signinvert = rs1_data[31] ^ rs2_data[31];
            mul_valid = !mul_ready;
            mul_factor0 = rs1_data[31] ? -rs1_data : rs1_data;
            mul_factor1 = rs2_data[31] ? -rs2_data : rs2_data;
            if(mul_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_MULH;
            end
        end
        is_mulhu: begin
            e2f_ready = 0;
            mul_signinvert = 0;
            mul_valid = !mul_ready;
            mul_factor0 = rs1_data;
            mul_factor1 = rs2_data;
            if(mul_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_MULH;
            end
        end
        is_mulhsu: begin
            e2f_ready = 0;
            mul_signinvert = rs1_data[31];
            mul_valid = !mul_ready;
            mul_factor0 = rs1_data[31] ? -rs1_data : rs1_data;
            mul_factor1 = rs2_data;
            if(mul_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_MULH;
            end
        end
        is_divu: begin
            e2f_ready = 0;
            div_fetch = !div_ready;
            div_signinvert = 0;
            div_dividend = rs1_data;
            div_divisor = rs2_data;
            // TODO: Division by zero
            if(div_ready && div_division_by_zero) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_MINUS_ONE;
            end else if(div_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_DIV;
            end
        end
        is_div: begin
            e2f_ready = 0;
            div_fetch = !div_ready;
            div_signinvert = rs1_data[31] ^ rs2_data[31];
            div_dividend = rs1_data[31] ? -rs1_data : rs1_data;
            div_divisor = rs2_data[31] ? -rs2_data : rs2_data;
            // TODO: Division by zero
            if(div_ready && div_division_by_zero) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_MINUS_ONE;
            end else if(div_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_DIV;
            end
        end
        is_remu: begin
            e2f_ready = 0;
            div_fetch = !div_ready;
            div_signinvert = 0;
            div_dividend = rs1_data;
            div_divisor = rs2_data;
            if(div_ready && div_division_by_zero) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_RS1;
            end else if(div_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_REM;
            end
        end
        is_rem: begin
            e2f_ready = 0;
            div_fetch = !div_ready;
            div_signinvert = rs1_data[31];
            div_dividend = rs1_data[31] ? -rs1_data : rs1_data;
            div_divisor = rs2_data[31] ? -rs2_data : rs2_data;
            if(div_ready && div_division_by_zero) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_RS1;
            end else if(div_ready) begin
                e2f_ready = 1;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_REM;
            end
        end
        is_op_imm, is_op: begin
            rd_write = (rd_addr != 0);
            rd_sel = `RD_ALU;
            illegal_instruction = alu_illegal_instruction;
            e2f_ready = 1;
        end
        is_jal: begin
            e2f_branchtaken = 1;
            e2f_branchtarget = f2e_pc + immgen_jal_offset;
            rd_write = (rd_addr != 0);
            rd_sel = `RD_PC_PLUS_4;
            e2f_ready = 1;
        end
        is_jalr: begin
            e2f_ready = 1;
            if(funct3 != 0) begin
                illegal_instruction = 1;
            end else begin
                e2f_branchtaken = 1;
                e2f_branchtarget = rs1_data + immgen_simm12;
                rd_write = (rd_addr != 0);
                rd_sel = `RD_PC_PLUS_4;
            end
        end
        is_branch: begin
            e2f_ready = 1;
            if(brcond_illegal_instruction) begin
                illegal_instruction = 1;
            end else begin
                e2f_branchtaken = brcond_branchtaken;
                e2f_branchtarget = f2e_pc + immgen_branch_offset;
            end
        end
        is_lui: begin
            e2f_ready = 1;
            rd_write = (rd_addr != 0);
            rd_sel = `RD_LUI;
        end
        is_auipc: begin
            e2f_ready = 1;
            rd_write = (rd_addr != 0);
            rd_sel = `RD_AUIPC;
        end
        is_load: begin
            e2f_ready = 0;
            c_address = rs1_data + immgen_simm12;
            c_cmd = `CACHE_CMD_LOAD;
            if(!dcache_command_issued) begin
                
            end else begin
                if(dcache_response_done) begin
                    rd_sel = `RD_DCACHE;
                    rd_write = (rd_addr != 0);
                    c_cmd = `CACHE_CMD_NONE;
                    e2f_ready = 1;
                end else if(dcache_response_error) begin
                    dcache_exc = 1;
                    e2f_ready = 1;
                    c_cmd = `CACHE_CMD_NONE;
                    if(c_response == `CACHE_RESPONSE_MISSALIGNED)
                        dcache_exc_cause = `EXCEPTION_CODE_LOAD_ADDRESS_MISALIGNED;
                    else if(c_response == `CACHE_RESPONSE_PAGEFAULT)
                        dcache_exc_cause = `EXCEPTION_CODE_LOAD_PAGE_FAULT;
                    else if(c_response == `CACHE_RESPONSE_ACCESSFAULT)
                        dcache_exc_cause = `EXCEPTION_CODE_LOAD_ACCESS_FAULT;
                end
            end
        end
        is_store: begin
            c_address = rs1_data + immgen_store_offset;
            c_cmd = `CACHE_CMD_STORE;
            if(funct3[2] != 0) begin
                c_cmd = `CACHE_CMD_NONE;
                illegal_instruction = 1;
                e2f_ready = 1;
            end else if(!dcache_command_issued) begin
                c_cmd = `CACHE_CMD_STORE;
                e2f_ready = 0;
            end else if(dcache_command_issued) begin
                e2f_ready = 0;
                c_cmd = `CACHE_CMD_STORE;
                if(dcache_response_done) begin
                    e2f_ready = 1;
                    c_cmd = `CACHE_CMD_NONE;
                end else if(dcache_response_error) begin
                    dcache_exc = 1;
                    e2f_ready = 1;
                    c_cmd = `CACHE_CMD_NONE;
                    if(c_response == `CACHE_RESPONSE_MISSALIGNED)
                        dcache_exc_cause = `EXCEPTION_CODE_STORE_ADDRESS_MISALIGNED;
                    else if(c_response == `CACHE_RESPONSE_PAGEFAULT)
                        dcache_exc_cause = `EXCEPTION_CODE_STORE_PAGE_FAULT;
                    else if(c_response == `CACHE_RESPONSE_ACCESSFAULT)
                        dcache_exc_cause = `EXCEPTION_CODE_STORE_ACCESS_FAULT;
                end
            end
        end
        is_fence: begin
            // Not implemented, just yet
            if(f2e_instr[31:28] == 4'b0000) begin
                if(!dcache_command_issued) begin
                    c_cmd = `CACHE_CMD_FLUSH_ALL;
                    e2f_ready = 0;
                end else if(dcache_command_issued) begin
                    e2f_ready = 0;
                    c_cmd = `CACHE_CMD_FLUSH_ALL;
                    if(dcache_response_done) begin
                        e2f_flush = 1;
                        e2f_ready = 1;
                        c_cmd = `CACHE_CMD_NONE;
                    end
                end
            end else begin
                illegal_instruction = 1;
            end
        end
        is_system: begin
            //illegal_instruction = 1;
            if(is_ebreak) begin
                e2f_ready = 0;
                e2debug_machine_ebreak = 1;
            end
            // Just temporary thing, pause on ebreak, for testing purposes

            // Handle CSR but with 1 cycle delay

            // TODO: Handle EBREAK, ECALL
            if(is_ecall) begin
                e2f_cmd = `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN;

                csr_cmd = `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN;
                csr_exc_cause = `EXCEPTION_CODE_ILLEGAL_INSTRUCTION;
                if(csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_MACHINE)
                    csr_exc_cause = ;
                else if(csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_SUPERVISOR)
                    csr_exc_cause = ;
                else if
            end else if(is_ebreak) begin
                if(csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_MACHINE) begin
                    e2debug_machine_ebreak = 1;
                end
            end else if(is_wfi && !csr_mstatus_tw) begin
                
            end else if(is_mret && (csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_MACHINE)) begin

            end else if(is_sret && !csr_mstatus_tsr && ((csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_MACHINE) || (csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_SUPERVISOR))) begin
                
            end else begin
                illegal_instruction = 1;
            end
        end
        default: begin
            illegal_instruction = 1;
        end
    endcase

    // TODO: Check csr_exc_privilege
    if(illegal_instruction) begin
        e2f_ready = 1;
        e2f_cmd = `ARMLEOCPU_E2F_CMD_BUBBLE_BRANCH;
        // e2f_bubble_exc_start_target = csr_next_pc;
        csr_cmd = `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN;
        csr_exc_cause = `EXCEPTION_CODE_ILLEGAL_INSTRUCTION;

    end else if(dcache_exc) begin
        e2f_ready = 1;
        e2f_cmd = `ARMLEOCPU_E2F_CMD_BUBBLE_BRANCH;

        csr_cmd = `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN;
        csr_exc_cause = dcache_exc_cause;
    end
    
    csr_exc_epc = f2e_epc;
    csr_exc_cause = f2e_cause;
    if(csr_mcurrent_privilege == `ARMLEOCPU_PRIVILEGE_MACHINE)
        csr_exc_privilege = `ARMLEOCPU_PRIVILEGE_MACHINE;
    else
        csr_exc_privilege = csr_medeleg[f2e_cause & ~] ? `ARMLEOCPU_PRIVILEGE_SUPERVISOR : `ARMLEOCPU_PRIVILEGE_MACHINE;
    if(f2e_exc_start) begin
        // TODO: ASSERT f2e_instr == NOP
        e2f_ready = 1;
        csr_exc_cmd = `ARMLEOCPU_CSR_CMD_INTERRUPT_BEGIN;
    end else if(f2e_exc_return) begin
        = ;
    end
end

always @(posedge clk) begin
    if(!rst_n) begin
        dcache_command_issued <= 0;
        csr_done <= 0;
    end else if(c_reset_done) begin
        if(illegal_instruction) begin
            `ifdef DEBUG_EXECUTE
                $display("[%m][%d][Execute] Illegal instruction, f2e_instr = 0x%X, f2e_pc = 0x%X", $time, f2e_instr, f2e_pc);
            `endif
        end else begin
            if(is_mulhu || is_mul || is_mulh || is_mulhsu) begin
                
                if(mul_ready) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] MUL instruction, done, f2e_instr = 0x%X, f2e_pc = 0x%X, rs1_data = 0x%X, rs2_data = 0x%X, rd_wdata = 0x%X, rd_write = %d", $time, f2e_instr, f2e_pc, rs1_data, rs2_data, rd_wdata, rd_write);
                    `endif
                end
            end else if(is_div || is_divu) begin
                if(div_ready) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] DIV instruction, done, f2e_instr = 0x%X, f2e_pc = 0x%X, rs1_data = 0x%X, rs2_data = 0x%X, rd_wdata = 0x%X, rd_write = %d", $time, f2e_instr, f2e_pc, rs1_data, rs2_data, rd_wdata, rd_write);
                    `endif
                end
            end else if(is_rem || is_remu) begin
                if(div_ready) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] REM instruction, done, f2e_instr = 0x%X, f2e_pc = 0x%X, rs1_data = 0x%X, rs2_data = 0x%X, rd_wdata = 0x%X, rd_write = %d", $time, f2e_instr, f2e_pc, rs1_data, rs2_data, rd_wdata, rd_write);
                    `endif
                end
            end else if(is_op || is_op_imm) begin
                if(alu_illegal_instruction) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] ALU Illegal instruction, f2e_instr = 0x%X, f2e_pc = 0x%X", $time, f2e_instr, f2e_pc);
                    `endif
                end
                if(is_op) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] ALU instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, rs1_data = 0x%X, rs2_data = 0x%X, rd_wdata = 0x%X, rd_write = %d", $time, f2e_instr, f2e_pc, rs1_data, rs2_data, rd_wdata, rd_write);
                    `endif
                end
                if(is_op_imm) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] ALU IMM instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, rs1_data = 0x%X, immgen_simm12 = 0x%X, rd_wdata = 0x%X, rd_write = %d", $time, f2e_instr, f2e_pc, rs1_data, immgen_simm12, rd_wdata, rd_write);
                    `endif
                end
            end else if(is_jal) begin
                `ifdef DEBUG_EXECUTE
                    $display("[%m][%d][Execute] JAL instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, e2f_branchtarget = 0x%X, immgen_jal_offset = 0x%X", $time, f2e_instr, f2e_pc, e2f_branchtarget, immgen_jal_offset);
                `endif
            end else if(is_jalr) begin
                `ifdef DEBUG_EXECUTE
                    $display("[%m][%d][Execute] JALR instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, e2f_branchtarget = 0x%X", $time, f2e_instr, f2e_pc, e2f_branchtarget);
                `endif
            end else if(is_branch) begin
                if(e2f_branchtaken) begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] Branch taken, f2e_instr = 0x%X, f2e_pc = 0x%X, e2f_branchtarget = 0x%X, rs1_data = 0x%X, rs2_data = 0x%X", $time, f2e_instr, f2e_pc, e2f_branchtarget, rs1_data, rs2_data);
                    `endif
                end else begin
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] Branch not taken, f2e_instr = 0x%X, f2e_pc = 0x%X", $time, f2e_instr, f2e_pc);
                    `endif
                end
            end else if(is_lui) begin
                `ifdef DEBUG_EXECUTE
                    $display("[%m][%d][Execute] LUI instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, rd_wdata = 0x%X", $time, f2e_instr, f2e_pc, rd_wdata);
                `endif
            end else if(is_auipc) begin
                `ifdef DEBUG_EXECUTE
                    $display("[%m][%d][Execute] AUIPC instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, rd_wdata = 0x%X", $time, f2e_instr, f2e_pc, rd_wdata);
                `endif
            end else if(is_load) begin
                if(!dcache_command_issued) begin
                    dcache_command_issued <= 1;
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] Load instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, c_response = , c_load_type = ,", $time, f2e_instr, f2e_pc);
                    `endif
                end else begin
                    if(dcache_response_done) begin
                        `ifdef DEBUG_EXECUTE
                            $display("[%m][%d][Execute] Load instruction, done, f2e_instr = 0x%X, f2e_pc = 0x%X, c_address = 0x%X, c_response = 0x%X, c_load_type = 0x%X, c_load_data = 0x%X", $time, f2e_instr, f2e_pc, c_address, c_response, c_load_type, c_load_data);
                        `endif
                        dcache_command_issued <= 0;
                    end else if(dcache_response_error) begin
                        `ifdef DEBUG_EXECUTE
                            $display("[%m][%d][Execute] Load instruction, error, f2e_instr = 0x%X, f2e_pc = 0x%X, c_address = 0x%X, c_response = 0x%X, c_load_type = 0x%X", $time, f2e_instr, f2e_pc, c_address, c_response, c_load_type);
                        `endif
                        dcache_command_issued <= 0;
                    end
                end
            end else if(is_store) begin
                if(!dcache_command_issued) begin
                    dcache_command_issued <= 1;
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] Store instruction, f2e_instr = 0x%X, f2e_pc = 0x%X, c_store_type = 0x%X", $time, f2e_instr, f2e_pc, c_store_type);
                    `endif
                end else begin
                    if(dcache_response_done) begin
                        `ifdef DEBUG_EXECUTE
                            $display("[%m][%d][Execute]  Store instruction, done, f2e_instr = 0x%X, f2e_pc = 0x%X, c_address = 0x%X, c_response = 0x%X, c_store_type = 0x%X, c_store_data = 0x%X", $time, f2e_instr, f2e_pc, c_address, c_response, c_store_type, c_store_data);
                        `endif
                        dcache_command_issued <= 0;
                    end else if(dcache_response_error) begin
                        dcache_command_issued <= 0;
                        `ifdef DEBUG_EXECUTE
                            $display("[%m][%d][Execute] Store instruction, error, f2e_instr = 0x%X, f2e_pc = 0x%X, c_address = 0x%X, c_response = 0x%X, c_load_type = 0x%X", $time, f2e_instr, f2e_pc, c_address, c_response, c_store_type);
                        `endif
                    end
                end
            end else if(is_fence) begin
                if(!dcache_command_issued) begin
                    dcache_command_issued <= 1'b1;
                    `ifdef DEBUG_EXECUTE
                        $display("[%m][%d][Execute] Fence instruction, f2e_instr = 0x%X, f2e_pc = 0x%X", $time, f2e_instr, f2e_pc);
                    `endif
                end else if(dcache_command_issued) begin
                    if(dcache_response_done) begin
                        dcache_command_issued <= 1'b0;
                        `ifdef DEBUG_EXECUTE
                            $display("[%m][%d][Execute] Fence instruction, done, f2e_instr = 0x%X, f2e_pc = 0x%X", $time, f2e_instr, f2e_pc);
                        `endif
                    end
                end
            end
        end
    end
end

endmodule