
localparam OPCODE_LUI    = 7'b0110111;
localparam OPCODE_AUIPC  = 7'b0010111;
localparam OPCODE_JAL    = 7'b1101111;
localparam OPCODE_JALR   = 7'b1100111;
localparam OPCODE_BRANCH = 7'b1100011;
localparam OPCODE_LOAD   = 7'b0000011;
localparam OPCODE_STORE  = 7'b0100011;
localparam OPCODE_ALUI   = 7'b0010011;
localparam OPCODE_ALU    = 7'b0110011;
localparam OPCODE_MISCMEM= 7'b0001111;
localparam OPCODE_SYSTEM = 7'b1110011;