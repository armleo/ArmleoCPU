module armleocpu_ptw(
    input clk,
    input async_rst_n,

    
);



endmodule