`define COREVX_PRIVILEGE_USER (2'b00)
`define COREVX_PRIVILEGE_SUPERVISOR (2'b01)
`define COREVX_PRIVILEGE_MACHINE (2'b11)