module armleocpu_execute (
    input clk,
    input rst_n,

    input [31:0] rs1_rdata,
    input [31:0] rs2_rdata,


    
    
);
    