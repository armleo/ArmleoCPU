
`undef ACCESS_PACKED
