/*
module armleocpu_decode (
// Fetch unit
    input      [31:0]       f2d_instr,
    input                   f2d_instr_valid,
    input      [31:0]       f2d_pc,
    input                   f2d_exc_start,
    input      [1:0]        f2d_exc_privilege,
    input      [31:0]       f2d_epc,
    input      [31:0]       f2d_cause,

    output reg              e2d_ready,
    output reg [`ARMLEOCPU_e2d_CMD_WIDTH-1:0]
                            e2d_cmd,
    output reg [31:0]       e2d_bubble_jump_target,
    output reg [31:0]       e2d_branchtarget,
);



endmodule*/
