`define TLB_CMD_NONE (2'b00)
`define TLB_CMD_RESOLVE (2'b01)
`define TLB_CMD_WRITE (2'b10)
`define TLB_CMD_INVALIDATE (2'b11)