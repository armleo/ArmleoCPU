
initial begin
	$dumpfile(`SIMRESULT);
	$dumpvars(0, `TOP);
end
