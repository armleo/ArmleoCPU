`define CSR_EXC_NONE (2'd0)
`define CSR_EXC_START (2'd1)
`define CSR_EXC_MRET (2'd2)
`define CSR_EXC_SRET (2'd3)

`define CSR_CMD_NONE (4'd0)
`define CSR_CMD_READ (4'd1)
`define CSR_CMD_WRITE (4'd2)
`define CSR_CMD_READ_WRITE (4'd3)
`define CSR_CMD_READ_SET (4'd4)
`define CSR_CMD_READ_CLEAR (4'd5)
`define CSR_CMD_MRET (4'd6)
`define CSR_CMD_SRET (4'd7)
`define CSR_CMD_INTERRUPT_BEGIN (4'd8)